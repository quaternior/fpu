// Wallace tree
module mult(
    output [47:0] product,
    input [23:0] A, B
);
    assign product = A * B;

endmodule
