// Wallace tree
module mult(
    output [47:0] product,
    input [23:0] A, B
);

wire [46:0] partial_products[23:0];

// i=1, j=23 => 1-(1+23-23)
// Partial product generation
genvar i, j;
generate
    for (i = 0; i < 24; i = i + 1) begin : pp_generation
        for (j = 0; j < 24; j = j + 1) begin : pp_gen
            if(i+j>23) begin  //If column idx is larger than bit width,
                assign partial_products[23-j][i+j] = A[j] & B[i];
            end
            else begin
                assign partial_products[i][i+j] = A[j] & B[i];
            end
        end
    end
endgenerate

// Final addition
// assign product = L7[22] + (carry[21] << 1);

wire [47:0] L1[22:0];
wire [47:0] L2[22:0];
wire [47:0] L3[22:0];
wire [47:0] L4[22:0];
wire [47:0] L5[22:0];
wire [47:0] L6[22:0];
wire [47:0] L7[22:0];

assign product[7:0] = L7[0][7:0];
//40-bit adder
adder adder_inst(product[47:8], L7[0][47:8], L7[1][47:8]);
wire [47:0] product_correct;
assign product_correct[7:0] = L7[0][7:0];
adder_correct adder_correct_inst(product_correct[47:8], L7[0][47:8], {1'b0, L7[1][46:8]});
//Auto-generated by python
assign L1[0][0] = partial_products[0][0];

ha ha_L1_0(L1[0][1], L1[0][1+1], partial_products[0][1], partial_products[0+1][1]);

fa fa_L1_1(L1[1][2], L1[0][2+1], partial_products[0][2], partial_products[0+1][2], partial_products[0+2][2]);

assign L1[1][3] = partial_products[0][3];
fa fa_L1_2(L1[2][3], L1[0][3+1], partial_products[1][3], partial_products[1+1][3], partial_products[1+2][3]);

ha ha_L1_3(L1[1][4], L1[0][4+1], partial_products[0][4], partial_products[0+1][4]);
fa fa_L1_4(L1[2][4], L1[1][4+1], partial_products[2][4], partial_products[2+1][4], partial_products[2+2][4]);

fa fa_L1_5(L1[2][5], L1[0][5+1], partial_products[0][5], partial_products[0+1][5], partial_products[0+2][5]);
fa fa_L1_6(L1[3][5], L1[1][5+1], partial_products[3][5], partial_products[3+1][5], partial_products[3+2][5]);

assign L1[2][6] = partial_products[0][6];
fa fa_L1_7(L1[3][6], L1[0][6+1], partial_products[1][6], partial_products[1+1][6], partial_products[1+2][6]);
fa fa_L1_8(L1[4][6], L1[1][6+1], partial_products[4][6], partial_products[4+1][6], partial_products[4+2][6]);

ha ha_L1_9(L1[2][7], L1[0][7+1], partial_products[0][7], partial_products[0+1][7]);
fa fa_L1_10(L1[3][7], L1[1][7+1], partial_products[2][7], partial_products[2+1][7], partial_products[2+2][7]);
fa fa_L1_11(L1[4][7], L1[2][7+1], partial_products[5][7], partial_products[5+1][7], partial_products[5+2][7]);

fa fa_L1_12(L1[3][8], L1[0][8+1], partial_products[0][8], partial_products[0+1][8], partial_products[0+2][8]);
fa fa_L1_13(L1[4][8], L1[1][8+1], partial_products[3][8], partial_products[3+1][8], partial_products[3+2][8]);
fa fa_L1_14(L1[5][8], L1[2][8+1], partial_products[6][8], partial_products[6+1][8], partial_products[6+2][8]);

assign L1[3][9] = partial_products[0][9];
fa fa_L1_15(L1[4][9], L1[0][9+1], partial_products[1][9], partial_products[1+1][9], partial_products[1+2][9]);
fa fa_L1_16(L1[5][9], L1[1][9+1], partial_products[4][9], partial_products[4+1][9], partial_products[4+2][9]);
fa fa_L1_17(L1[6][9], L1[2][9+1], partial_products[7][9], partial_products[7+1][9], partial_products[7+2][9]);

ha ha_L1_18(L1[3][10], L1[0][10+1], partial_products[0][10], partial_products[0+1][10]);
fa fa_L1_19(L1[4][10], L1[1][10+1], partial_products[2][10], partial_products[2+1][10], partial_products[2+2][10]);
fa fa_L1_20(L1[5][10], L1[2][10+1], partial_products[5][10], partial_products[5+1][10], partial_products[5+2][10]);
fa fa_L1_21(L1[6][10], L1[3][10+1], partial_products[8][10], partial_products[8+1][10], partial_products[8+2][10]);

fa fa_L1_22(L1[4][11], L1[0][11+1], partial_products[0][11], partial_products[0+1][11], partial_products[0+2][11]);
fa fa_L1_23(L1[5][11], L1[1][11+1], partial_products[3][11], partial_products[3+1][11], partial_products[3+2][11]);
fa fa_L1_24(L1[6][11], L1[2][11+1], partial_products[6][11], partial_products[6+1][11], partial_products[6+2][11]);
fa fa_L1_25(L1[7][11], L1[3][11+1], partial_products[9][11], partial_products[9+1][11], partial_products[9+2][11]);

assign L1[4][12] = partial_products[0][12];
fa fa_L1_26(L1[5][12], L1[0][12+1], partial_products[1][12], partial_products[1+1][12], partial_products[1+2][12]);
fa fa_L1_27(L1[6][12], L1[1][12+1], partial_products[4][12], partial_products[4+1][12], partial_products[4+2][12]);
fa fa_L1_28(L1[7][12], L1[2][12+1], partial_products[7][12], partial_products[7+1][12], partial_products[7+2][12]);
fa fa_L1_29(L1[8][12], L1[3][12+1], partial_products[10][12], partial_products[10+1][12], partial_products[10+2][12]);

ha ha_L1_30(L1[4][13], L1[0][13+1], partial_products[0][13], partial_products[0+1][13]);
fa fa_L1_31(L1[5][13], L1[1][13+1], partial_products[2][13], partial_products[2+1][13], partial_products[2+2][13]);
fa fa_L1_32(L1[6][13], L1[2][13+1], partial_products[5][13], partial_products[5+1][13], partial_products[5+2][13]);
fa fa_L1_33(L1[7][13], L1[3][13+1], partial_products[8][13], partial_products[8+1][13], partial_products[8+2][13]);
fa fa_L1_34(L1[8][13], L1[4][13+1], partial_products[11][13], partial_products[11+1][13], partial_products[11+2][13]);

fa fa_L1_35(L1[5][14], L1[0][14+1], partial_products[0][14], partial_products[0+1][14], partial_products[0+2][14]);
fa fa_L1_36(L1[6][14], L1[1][14+1], partial_products[3][14], partial_products[3+1][14], partial_products[3+2][14]);
fa fa_L1_37(L1[7][14], L1[2][14+1], partial_products[6][14], partial_products[6+1][14], partial_products[6+2][14]);
fa fa_L1_38(L1[8][14], L1[3][14+1], partial_products[9][14], partial_products[9+1][14], partial_products[9+2][14]);
fa fa_L1_39(L1[9][14], L1[4][14+1], partial_products[12][14], partial_products[12+1][14], partial_products[12+2][14]);

assign L1[5][15] = partial_products[0][15];
fa fa_L1_40(L1[6][15], L1[0][15+1], partial_products[1][15], partial_products[1+1][15], partial_products[1+2][15]);
fa fa_L1_41(L1[7][15], L1[1][15+1], partial_products[4][15], partial_products[4+1][15], partial_products[4+2][15]);
fa fa_L1_42(L1[8][15], L1[2][15+1], partial_products[7][15], partial_products[7+1][15], partial_products[7+2][15]);
fa fa_L1_43(L1[9][15], L1[3][15+1], partial_products[10][15], partial_products[10+1][15], partial_products[10+2][15]);
fa fa_L1_44(L1[10][15], L1[4][15+1], partial_products[13][15], partial_products[13+1][15], partial_products[13+2][15]);

ha ha_L1_45(L1[5][16], L1[0][16+1], partial_products[0][16], partial_products[0+1][16]);
fa fa_L1_46(L1[6][16], L1[1][16+1], partial_products[2][16], partial_products[2+1][16], partial_products[2+2][16]);
fa fa_L1_47(L1[7][16], L1[2][16+1], partial_products[5][16], partial_products[5+1][16], partial_products[5+2][16]);
fa fa_L1_48(L1[8][16], L1[3][16+1], partial_products[8][16], partial_products[8+1][16], partial_products[8+2][16]);
fa fa_L1_49(L1[9][16], L1[4][16+1], partial_products[11][16], partial_products[11+1][16], partial_products[11+2][16]);
fa fa_L1_50(L1[10][16], L1[5][16+1], partial_products[14][16], partial_products[14+1][16], partial_products[14+2][16]);

fa fa_L1_51(L1[6][17], L1[0][17+1], partial_products[0][17], partial_products[0+1][17], partial_products[0+2][17]);
fa fa_L1_52(L1[7][17], L1[1][17+1], partial_products[3][17], partial_products[3+1][17], partial_products[3+2][17]);
fa fa_L1_53(L1[8][17], L1[2][17+1], partial_products[6][17], partial_products[6+1][17], partial_products[6+2][17]);
fa fa_L1_54(L1[9][17], L1[3][17+1], partial_products[9][17], partial_products[9+1][17], partial_products[9+2][17]);
fa fa_L1_55(L1[10][17], L1[4][17+1], partial_products[12][17], partial_products[12+1][17], partial_products[12+2][17]);
fa fa_L1_56(L1[11][17], L1[5][17+1], partial_products[15][17], partial_products[15+1][17], partial_products[15+2][17]);

assign L1[6][18] = partial_products[0][18];
fa fa_L1_57(L1[7][18], L1[0][18+1], partial_products[1][18], partial_products[1+1][18], partial_products[1+2][18]);
fa fa_L1_58(L1[8][18], L1[1][18+1], partial_products[4][18], partial_products[4+1][18], partial_products[4+2][18]);
fa fa_L1_59(L1[9][18], L1[2][18+1], partial_products[7][18], partial_products[7+1][18], partial_products[7+2][18]);
fa fa_L1_60(L1[10][18], L1[3][18+1], partial_products[10][18], partial_products[10+1][18], partial_products[10+2][18]);
fa fa_L1_61(L1[11][18], L1[4][18+1], partial_products[13][18], partial_products[13+1][18], partial_products[13+2][18]);
fa fa_L1_62(L1[12][18], L1[5][18+1], partial_products[16][18], partial_products[16+1][18], partial_products[16+2][18]);

ha ha_L1_63(L1[6][19], L1[0][19+1], partial_products[0][19], partial_products[0+1][19]);
fa fa_L1_64(L1[7][19], L1[1][19+1], partial_products[2][19], partial_products[2+1][19], partial_products[2+2][19]);
fa fa_L1_65(L1[8][19], L1[2][19+1], partial_products[5][19], partial_products[5+1][19], partial_products[5+2][19]);
fa fa_L1_66(L1[9][19], L1[3][19+1], partial_products[8][19], partial_products[8+1][19], partial_products[8+2][19]);
fa fa_L1_67(L1[10][19], L1[4][19+1], partial_products[11][19], partial_products[11+1][19], partial_products[11+2][19]);
fa fa_L1_68(L1[11][19], L1[5][19+1], partial_products[14][19], partial_products[14+1][19], partial_products[14+2][19]);
fa fa_L1_69(L1[12][19], L1[6][19+1], partial_products[17][19], partial_products[17+1][19], partial_products[17+2][19]);

fa fa_L1_70(L1[7][20], L1[0][20+1], partial_products[0][20], partial_products[0+1][20], partial_products[0+2][20]);
fa fa_L1_71(L1[8][20], L1[1][20+1], partial_products[3][20], partial_products[3+1][20], partial_products[3+2][20]);
fa fa_L1_72(L1[9][20], L1[2][20+1], partial_products[6][20], partial_products[6+1][20], partial_products[6+2][20]);
fa fa_L1_73(L1[10][20], L1[3][20+1], partial_products[9][20], partial_products[9+1][20], partial_products[9+2][20]);
fa fa_L1_74(L1[11][20], L1[4][20+1], partial_products[12][20], partial_products[12+1][20], partial_products[12+2][20]);
fa fa_L1_75(L1[12][20], L1[5][20+1], partial_products[15][20], partial_products[15+1][20], partial_products[15+2][20]);
fa fa_L1_76(L1[13][20], L1[6][20+1], partial_products[18][20], partial_products[18+1][20], partial_products[18+2][20]);

assign L1[7][21] = partial_products[0][21];
fa fa_L1_77(L1[8][21], L1[0][21+1], partial_products[1][21], partial_products[1+1][21], partial_products[1+2][21]);
fa fa_L1_78(L1[9][21], L1[1][21+1], partial_products[4][21], partial_products[4+1][21], partial_products[4+2][21]);
fa fa_L1_79(L1[10][21], L1[2][21+1], partial_products[7][21], partial_products[7+1][21], partial_products[7+2][21]);
fa fa_L1_80(L1[11][21], L1[3][21+1], partial_products[10][21], partial_products[10+1][21], partial_products[10+2][21]);
fa fa_L1_81(L1[12][21], L1[4][21+1], partial_products[13][21], partial_products[13+1][21], partial_products[13+2][21]);
fa fa_L1_82(L1[13][21], L1[5][21+1], partial_products[16][21], partial_products[16+1][21], partial_products[16+2][21]);
fa fa_L1_83(L1[14][21], L1[6][21+1], partial_products[19][21], partial_products[19+1][21], partial_products[19+2][21]);

ha ha_L1_84(L1[7][22], L1[0][22+1], partial_products[0][22], partial_products[0+1][22]);
fa fa_L1_85(L1[8][22], L1[1][22+1], partial_products[2][22], partial_products[2+1][22], partial_products[2+2][22]);
fa fa_L1_86(L1[9][22], L1[2][22+1], partial_products[5][22], partial_products[5+1][22], partial_products[5+2][22]);
fa fa_L1_87(L1[10][22], L1[3][22+1], partial_products[8][22], partial_products[8+1][22], partial_products[8+2][22]);
fa fa_L1_88(L1[11][22], L1[4][22+1], partial_products[11][22], partial_products[11+1][22], partial_products[11+2][22]);
fa fa_L1_89(L1[12][22], L1[5][22+1], partial_products[14][22], partial_products[14+1][22], partial_products[14+2][22]);
fa fa_L1_90(L1[13][22], L1[6][22+1], partial_products[17][22], partial_products[17+1][22], partial_products[17+2][22]);
fa fa_L1_91(L1[14][22], L1[7][22+1], partial_products[20][22], partial_products[20+1][22], partial_products[20+2][22]);

fa fa_L1_92(L1[8][23], L1[0][23+1], partial_products[0][23], partial_products[0+1][23], partial_products[0+2][23]);
fa fa_L1_93(L1[9][23], L1[1][23+1], partial_products[3][23], partial_products[3+1][23], partial_products[3+2][23]);
fa fa_L1_94(L1[10][23], L1[2][23+1], partial_products[6][23], partial_products[6+1][23], partial_products[6+2][23]);
fa fa_L1_95(L1[11][23], L1[3][23+1], partial_products[9][23], partial_products[9+1][23], partial_products[9+2][23]);
fa fa_L1_96(L1[12][23], L1[4][23+1], partial_products[12][23], partial_products[12+1][23], partial_products[12+2][23]);
fa fa_L1_97(L1[13][23], L1[5][23+1], partial_products[15][23], partial_products[15+1][23], partial_products[15+2][23]);
fa fa_L1_98(L1[14][23], L1[6][23+1], partial_products[18][23], partial_products[18+1][23], partial_products[18+2][23]);
fa fa_L1_99(L1[15][23], L1[7][23+1], partial_products[21][23], partial_products[21+1][23], partial_products[21+2][23]);

ha ha_L1_100(L1[8][24], L1[0][24+1], partial_products[0][24], partial_products[0+1][24]);
fa fa_L1_101(L1[9][24], L1[1][24+1], partial_products[2][24], partial_products[2+1][24], partial_products[2+2][24]);
fa fa_L1_102(L1[10][24], L1[2][24+1], partial_products[5][24], partial_products[5+1][24], partial_products[5+2][24]);
fa fa_L1_103(L1[11][24], L1[3][24+1], partial_products[8][24], partial_products[8+1][24], partial_products[8+2][24]);
fa fa_L1_104(L1[12][24], L1[4][24+1], partial_products[11][24], partial_products[11+1][24], partial_products[11+2][24]);
fa fa_L1_105(L1[13][24], L1[5][24+1], partial_products[14][24], partial_products[14+1][24], partial_products[14+2][24]);
fa fa_L1_106(L1[14][24], L1[6][24+1], partial_products[17][24], partial_products[17+1][24], partial_products[17+2][24]);
fa fa_L1_107(L1[15][24], L1[7][24+1], partial_products[20][24], partial_products[20+1][24], partial_products[20+2][24]);

assign L1[8][25] = partial_products[0][25];
fa fa_L1_108(L1[9][25], L1[0][25+1], partial_products[1][25], partial_products[1+1][25], partial_products[1+2][25]);
fa fa_L1_109(L1[10][25], L1[1][25+1], partial_products[4][25], partial_products[4+1][25], partial_products[4+2][25]);
fa fa_L1_110(L1[11][25], L1[2][25+1], partial_products[7][25], partial_products[7+1][25], partial_products[7+2][25]);
fa fa_L1_111(L1[12][25], L1[3][25+1], partial_products[10][25], partial_products[10+1][25], partial_products[10+2][25]);
fa fa_L1_112(L1[13][25], L1[4][25+1], partial_products[13][25], partial_products[13+1][25], partial_products[13+2][25]);
fa fa_L1_113(L1[14][25], L1[5][25+1], partial_products[16][25], partial_products[16+1][25], partial_products[16+2][25]);
fa fa_L1_114(L1[15][25], L1[6][25+1], partial_products[19][25], partial_products[19+1][25], partial_products[19+2][25]);

fa fa_L1_115(L1[7][26], L1[0][26+1], partial_products[0][26], partial_products[0+1][26], partial_products[0+2][26]);
fa fa_L1_116(L1[8][26], L1[1][26+1], partial_products[3][26], partial_products[3+1][26], partial_products[3+2][26]);
fa fa_L1_117(L1[9][26], L1[2][26+1], partial_products[6][26], partial_products[6+1][26], partial_products[6+2][26]);
fa fa_L1_118(L1[10][26], L1[3][26+1], partial_products[9][26], partial_products[9+1][26], partial_products[9+2][26]);
fa fa_L1_119(L1[11][26], L1[4][26+1], partial_products[12][26], partial_products[12+1][26], partial_products[12+2][26]);
fa fa_L1_120(L1[12][26], L1[5][26+1], partial_products[15][26], partial_products[15+1][26], partial_products[15+2][26]);
fa fa_L1_121(L1[13][26], L1[6][26+1], partial_products[18][26], partial_products[18+1][26], partial_products[18+2][26]);

ha ha_L1_122(L1[7][27], L1[0][27+1], partial_products[0][27], partial_products[0+1][27]);
fa fa_L1_123(L1[8][27], L1[1][27+1], partial_products[2][27], partial_products[2+1][27], partial_products[2+2][27]);
fa fa_L1_124(L1[9][27], L1[2][27+1], partial_products[5][27], partial_products[5+1][27], partial_products[5+2][27]);
fa fa_L1_125(L1[10][27], L1[3][27+1], partial_products[8][27], partial_products[8+1][27], partial_products[8+2][27]);
fa fa_L1_126(L1[11][27], L1[4][27+1], partial_products[11][27], partial_products[11+1][27], partial_products[11+2][27]);
fa fa_L1_127(L1[12][27], L1[5][27+1], partial_products[14][27], partial_products[14+1][27], partial_products[14+2][27]);
fa fa_L1_128(L1[13][27], L1[6][27+1], partial_products[17][27], partial_products[17+1][27], partial_products[17+2][27]);

assign L1[7][28] = partial_products[0][28];
fa fa_L1_129(L1[8][28], L1[0][28+1], partial_products[1][28], partial_products[1+1][28], partial_products[1+2][28]);
fa fa_L1_130(L1[9][28], L1[1][28+1], partial_products[4][28], partial_products[4+1][28], partial_products[4+2][28]);
fa fa_L1_131(L1[10][28], L1[2][28+1], partial_products[7][28], partial_products[7+1][28], partial_products[7+2][28]);
fa fa_L1_132(L1[11][28], L1[3][28+1], partial_products[10][28], partial_products[10+1][28], partial_products[10+2][28]);
fa fa_L1_133(L1[12][28], L1[4][28+1], partial_products[13][28], partial_products[13+1][28], partial_products[13+2][28]);
fa fa_L1_134(L1[13][28], L1[5][28+1], partial_products[16][28], partial_products[16+1][28], partial_products[16+2][28]);

fa fa_L1_135(L1[6][29], L1[0][29+1], partial_products[0][29], partial_products[0+1][29], partial_products[0+2][29]);
fa fa_L1_136(L1[7][29], L1[1][29+1], partial_products[3][29], partial_products[3+1][29], partial_products[3+2][29]);
fa fa_L1_137(L1[8][29], L1[2][29+1], partial_products[6][29], partial_products[6+1][29], partial_products[6+2][29]);
fa fa_L1_138(L1[9][29], L1[3][29+1], partial_products[9][29], partial_products[9+1][29], partial_products[9+2][29]);
fa fa_L1_139(L1[10][29], L1[4][29+1], partial_products[12][29], partial_products[12+1][29], partial_products[12+2][29]);
fa fa_L1_140(L1[11][29], L1[5][29+1], partial_products[15][29], partial_products[15+1][29], partial_products[15+2][29]);

ha ha_L1_141(L1[6][30], L1[0][30+1], partial_products[0][30], partial_products[0+1][30]);
fa fa_L1_142(L1[7][30], L1[1][30+1], partial_products[2][30], partial_products[2+1][30], partial_products[2+2][30]);
fa fa_L1_143(L1[8][30], L1[2][30+1], partial_products[5][30], partial_products[5+1][30], partial_products[5+2][30]);
fa fa_L1_144(L1[9][30], L1[3][30+1], partial_products[8][30], partial_products[8+1][30], partial_products[8+2][30]);
fa fa_L1_145(L1[10][30], L1[4][30+1], partial_products[11][30], partial_products[11+1][30], partial_products[11+2][30]);
fa fa_L1_146(L1[11][30], L1[5][30+1], partial_products[14][30], partial_products[14+1][30], partial_products[14+2][30]);

assign L1[6][31] = partial_products[0][31];
fa fa_L1_147(L1[7][31], L1[0][31+1], partial_products[1][31], partial_products[1+1][31], partial_products[1+2][31]);
fa fa_L1_148(L1[8][31], L1[1][31+1], partial_products[4][31], partial_products[4+1][31], partial_products[4+2][31]);
fa fa_L1_149(L1[9][31], L1[2][31+1], partial_products[7][31], partial_products[7+1][31], partial_products[7+2][31]);
fa fa_L1_150(L1[10][31], L1[3][31+1], partial_products[10][31], partial_products[10+1][31], partial_products[10+2][31]);
fa fa_L1_151(L1[11][31], L1[4][31+1], partial_products[13][31], partial_products[13+1][31], partial_products[13+2][31]);

fa fa_L1_152(L1[5][32], L1[0][32+1], partial_products[0][32], partial_products[0+1][32], partial_products[0+2][32]);
fa fa_L1_153(L1[6][32], L1[1][32+1], partial_products[3][32], partial_products[3+1][32], partial_products[3+2][32]);
fa fa_L1_154(L1[7][32], L1[2][32+1], partial_products[6][32], partial_products[6+1][32], partial_products[6+2][32]);
fa fa_L1_155(L1[8][32], L1[3][32+1], partial_products[9][32], partial_products[9+1][32], partial_products[9+2][32]);
fa fa_L1_156(L1[9][32], L1[4][32+1], partial_products[12][32], partial_products[12+1][32], partial_products[12+2][32]);

ha ha_L1_157(L1[5][33], L1[0][33+1], partial_products[0][33], partial_products[0+1][33]);
fa fa_L1_158(L1[6][33], L1[1][33+1], partial_products[2][33], partial_products[2+1][33], partial_products[2+2][33]);
fa fa_L1_159(L1[7][33], L1[2][33+1], partial_products[5][33], partial_products[5+1][33], partial_products[5+2][33]);
fa fa_L1_160(L1[8][33], L1[3][33+1], partial_products[8][33], partial_products[8+1][33], partial_products[8+2][33]);
fa fa_L1_161(L1[9][33], L1[4][33+1], partial_products[11][33], partial_products[11+1][33], partial_products[11+2][33]);

assign L1[5][34] = partial_products[0][34];
fa fa_L1_162(L1[6][34], L1[0][34+1], partial_products[1][34], partial_products[1+1][34], partial_products[1+2][34]);
fa fa_L1_163(L1[7][34], L1[1][34+1], partial_products[4][34], partial_products[4+1][34], partial_products[4+2][34]);
fa fa_L1_164(L1[8][34], L1[2][34+1], partial_products[7][34], partial_products[7+1][34], partial_products[7+2][34]);
fa fa_L1_165(L1[9][34], L1[3][34+1], partial_products[10][34], partial_products[10+1][34], partial_products[10+2][34]);

fa fa_L1_166(L1[4][35], L1[0][35+1], partial_products[0][35], partial_products[0+1][35], partial_products[0+2][35]);
fa fa_L1_167(L1[5][35], L1[1][35+1], partial_products[3][35], partial_products[3+1][35], partial_products[3+2][35]);
fa fa_L1_168(L1[6][35], L1[2][35+1], partial_products[6][35], partial_products[6+1][35], partial_products[6+2][35]);
fa fa_L1_169(L1[7][35], L1[3][35+1], partial_products[9][35], partial_products[9+1][35], partial_products[9+2][35]);

ha ha_L1_170(L1[4][36], L1[0][36+1], partial_products[0][36], partial_products[0+1][36]);
fa fa_L1_171(L1[5][36], L1[1][36+1], partial_products[2][36], partial_products[2+1][36], partial_products[2+2][36]);
fa fa_L1_172(L1[6][36], L1[2][36+1], partial_products[5][36], partial_products[5+1][36], partial_products[5+2][36]);
fa fa_L1_173(L1[7][36], L1[3][36+1], partial_products[8][36], partial_products[8+1][36], partial_products[8+2][36]);

assign L1[4][37] = partial_products[0][37];
fa fa_L1_174(L1[5][37], L1[0][37+1], partial_products[1][37], partial_products[1+1][37], partial_products[1+2][37]);
fa fa_L1_175(L1[6][37], L1[1][37+1], partial_products[4][37], partial_products[4+1][37], partial_products[4+2][37]);
fa fa_L1_176(L1[7][37], L1[2][37+1], partial_products[7][37], partial_products[7+1][37], partial_products[7+2][37]);

fa fa_L1_177(L1[3][38], L1[0][38+1], partial_products[0][38], partial_products[0+1][38], partial_products[0+2][38]);
fa fa_L1_178(L1[4][38], L1[1][38+1], partial_products[3][38], partial_products[3+1][38], partial_products[3+2][38]);
fa fa_L1_179(L1[5][38], L1[2][38+1], partial_products[6][38], partial_products[6+1][38], partial_products[6+2][38]);

ha ha_L1_180(L1[3][39], L1[0][39+1], partial_products[0][39], partial_products[0+1][39]);
fa fa_L1_181(L1[4][39], L1[1][39+1], partial_products[2][39], partial_products[2+1][39], partial_products[2+2][39]);
fa fa_L1_182(L1[5][39], L1[2][39+1], partial_products[5][39], partial_products[5+1][39], partial_products[5+2][39]);

assign L1[3][40] = partial_products[0][40];
fa fa_L1_183(L1[4][40], L1[0][40+1], partial_products[1][40], partial_products[1+1][40], partial_products[1+2][40]);
fa fa_L1_184(L1[5][40], L1[1][40+1], partial_products[4][40], partial_products[4+1][40], partial_products[4+2][40]);

fa fa_L1_185(L1[2][41], L1[0][41+1], partial_products[0][41], partial_products[0+1][41], partial_products[0+2][41]);
fa fa_L1_186(L1[3][41], L1[1][41+1], partial_products[3][41], partial_products[3+1][41], partial_products[3+2][41]);

ha ha_L1_187(L1[2][42], L1[0][42+1], partial_products[0][42], partial_products[0+1][42]);
fa fa_L1_188(L1[3][42], L1[1][42+1], partial_products[2][42], partial_products[2+1][42], partial_products[2+2][42]);

assign L1[2][43] = partial_products[0][43];
fa fa_L1_189(L1[3][43], L1[0][43+1], partial_products[1][43], partial_products[1+1][43], partial_products[1+2][43]);

fa fa_L1_190(L1[1][44], L1[0][44+1], partial_products[0][44], partial_products[0+1][44], partial_products[0+2][44]);

assign L1[1][45] = partial_products[0][45];
assign L1[2][45] = partial_products[1][45];

assign L1[0][46] = partial_products[0][46];


assign L2[0][0] = L1[0][0];

assign L2[0][1] = L1[0][1];

ha ha_L2_0(L2[0][2], L2[0][2+1], L1[0][2], L1[0+1][2]);

fa fa_L2_1(L2[1][3], L2[0][3+1], L1[0][3], L1[0+1][3], L1[0+2][3]);

fa fa_L2_2(L2[1][4], L2[0][4+1], L1[0][4], L1[0+1][4], L1[0+2][4]);

assign L2[1][5] = L1[0][5];
fa fa_L2_3(L2[2][5], L2[0][5+1], L1[1][5], L1[1+1][5], L1[1+2][5]);

ha ha_L2_4(L2[1][6], L2[0][6+1], L1[0][6], L1[0+1][6]);
fa fa_L2_5(L2[2][6], L2[1][6+1], L1[2][6], L1[2+1][6], L1[2+2][6]);

ha ha_L2_6(L2[2][7], L2[0][7+1], L1[0][7], L1[0+1][7]);
fa fa_L2_7(L2[3][7], L2[1][7+1], L1[2][7], L1[2+1][7], L1[2+2][7]);

fa fa_L2_8(L2[2][8], L2[0][8+1], L1[0][8], L1[0+1][8], L1[0+2][8]);
fa fa_L2_9(L2[3][8], L2[1][8+1], L1[3][8], L1[3+1][8], L1[3+2][8]);

assign L2[2][9] = L1[0][9];
fa fa_L2_10(L2[3][9], L2[0][9+1], L1[1][9], L1[1+1][9], L1[1+2][9]);
fa fa_L2_11(L2[4][9], L2[1][9+1], L1[4][9], L1[4+1][9], L1[4+2][9]);

assign L2[2][10] = L1[0][10];
fa fa_L2_12(L2[3][10], L2[0][10+1], L1[1][10], L1[1+1][10], L1[1+2][10]);
fa fa_L2_13(L2[4][10], L2[1][10+1], L1[4][10], L1[4+1][10], L1[4+2][10]);

ha ha_L2_14(L2[2][11], L2[0][11+1], L1[0][11], L1[0+1][11]);
fa fa_L2_15(L2[3][11], L2[1][11+1], L1[2][11], L1[2+1][11], L1[2+2][11]);
fa fa_L2_16(L2[4][11], L2[2][11+1], L1[5][11], L1[5+1][11], L1[5+2][11]);

fa fa_L2_17(L2[3][12], L2[0][12+1], L1[0][12], L1[0+1][12], L1[0+2][12]);
fa fa_L2_18(L2[4][12], L2[1][12+1], L1[3][12], L1[3+1][12], L1[3+2][12]);
fa fa_L2_19(L2[5][12], L2[2][12+1], L1[6][12], L1[6+1][12], L1[6+2][12]);

fa fa_L2_20(L2[3][13], L2[0][13+1], L1[0][13], L1[0+1][13], L1[0+2][13]);
fa fa_L2_21(L2[4][13], L2[1][13+1], L1[3][13], L1[3+1][13], L1[3+2][13]);
fa fa_L2_22(L2[5][13], L2[2][13+1], L1[6][13], L1[6+1][13], L1[6+2][13]);

assign L2[3][14] = L1[0][14];
fa fa_L2_23(L2[4][14], L2[0][14+1], L1[1][14], L1[1+1][14], L1[1+2][14]);
fa fa_L2_24(L2[5][14], L2[1][14+1], L1[4][14], L1[4+1][14], L1[4+2][14]);
fa fa_L2_25(L2[6][14], L2[2][14+1], L1[7][14], L1[7+1][14], L1[7+2][14]);

ha ha_L2_26(L2[3][15], L2[0][15+1], L1[0][15], L1[0+1][15]);
fa fa_L2_27(L2[4][15], L2[1][15+1], L1[2][15], L1[2+1][15], L1[2+2][15]);
fa fa_L2_28(L2[5][15], L2[2][15+1], L1[5][15], L1[5+1][15], L1[5+2][15]);
fa fa_L2_29(L2[6][15], L2[3][15+1], L1[8][15], L1[8+1][15], L1[8+2][15]);

ha ha_L2_30(L2[4][16], L2[0][16+1], L1[0][16], L1[0+1][16]);
fa fa_L2_31(L2[5][16], L2[1][16+1], L1[2][16], L1[2+1][16], L1[2+2][16]);
fa fa_L2_32(L2[6][16], L2[2][16+1], L1[5][16], L1[5+1][16], L1[5+2][16]);
fa fa_L2_33(L2[7][16], L2[3][16+1], L1[8][16], L1[8+1][16], L1[8+2][16]);

fa fa_L2_34(L2[4][17], L2[0][17+1], L1[0][17], L1[0+1][17], L1[0+2][17]);
fa fa_L2_35(L2[5][17], L2[1][17+1], L1[3][17], L1[3+1][17], L1[3+2][17]);
fa fa_L2_36(L2[6][17], L2[2][17+1], L1[6][17], L1[6+1][17], L1[6+2][17]);
fa fa_L2_37(L2[7][17], L2[3][17+1], L1[9][17], L1[9+1][17], L1[9+2][17]);

assign L2[4][18] = L1[0][18];
fa fa_L2_38(L2[5][18], L2[0][18+1], L1[1][18], L1[1+1][18], L1[1+2][18]);
fa fa_L2_39(L2[6][18], L2[1][18+1], L1[4][18], L1[4+1][18], L1[4+2][18]);
fa fa_L2_40(L2[7][18], L2[2][18+1], L1[7][18], L1[7+1][18], L1[7+2][18]);
fa fa_L2_41(L2[8][18], L2[3][18+1], L1[10][18], L1[10+1][18], L1[10+2][18]);

assign L2[4][19] = L1[0][19];
fa fa_L2_42(L2[5][19], L2[0][19+1], L1[1][19], L1[1+1][19], L1[1+2][19]);
fa fa_L2_43(L2[6][19], L2[1][19+1], L1[4][19], L1[4+1][19], L1[4+2][19]);
fa fa_L2_44(L2[7][19], L2[2][19+1], L1[7][19], L1[7+1][19], L1[7+2][19]);
fa fa_L2_45(L2[8][19], L2[3][19+1], L1[10][19], L1[10+1][19], L1[10+2][19]);

ha ha_L2_46(L2[4][20], L2[0][20+1], L1[0][20], L1[0+1][20]);
fa fa_L2_47(L2[5][20], L2[1][20+1], L1[2][20], L1[2+1][20], L1[2+2][20]);
fa fa_L2_48(L2[6][20], L2[2][20+1], L1[5][20], L1[5+1][20], L1[5+2][20]);
fa fa_L2_49(L2[7][20], L2[3][20+1], L1[8][20], L1[8+1][20], L1[8+2][20]);
fa fa_L2_50(L2[8][20], L2[4][20+1], L1[11][20], L1[11+1][20], L1[11+2][20]);

fa fa_L2_51(L2[5][21], L2[0][21+1], L1[0][21], L1[0+1][21], L1[0+2][21]);
fa fa_L2_52(L2[6][21], L2[1][21+1], L1[3][21], L1[3+1][21], L1[3+2][21]);
fa fa_L2_53(L2[7][21], L2[2][21+1], L1[6][21], L1[6+1][21], L1[6+2][21]);
fa fa_L2_54(L2[8][21], L2[3][21+1], L1[9][21], L1[9+1][21], L1[9+2][21]);
fa fa_L2_55(L2[9][21], L2[4][21+1], L1[12][21], L1[12+1][21], L1[12+2][21]);

fa fa_L2_56(L2[5][22], L2[0][22+1], L1[0][22], L1[0+1][22], L1[0+2][22]);
fa fa_L2_57(L2[6][22], L2[1][22+1], L1[3][22], L1[3+1][22], L1[3+2][22]);
fa fa_L2_58(L2[7][22], L2[2][22+1], L1[6][22], L1[6+1][22], L1[6+2][22]);
fa fa_L2_59(L2[8][22], L2[3][22+1], L1[9][22], L1[9+1][22], L1[9+2][22]);
fa fa_L2_60(L2[9][22], L2[4][22+1], L1[12][22], L1[12+1][22], L1[12+2][22]);

assign L2[5][23] = L1[0][23];
fa fa_L2_61(L2[6][23], L2[0][23+1], L1[1][23], L1[1+1][23], L1[1+2][23]);
fa fa_L2_62(L2[7][23], L2[1][23+1], L1[4][23], L1[4+1][23], L1[4+2][23]);
fa fa_L2_63(L2[8][23], L2[2][23+1], L1[7][23], L1[7+1][23], L1[7+2][23]);
fa fa_L2_64(L2[9][23], L2[3][23+1], L1[10][23], L1[10+1][23], L1[10+2][23]);
fa fa_L2_65(L2[10][23], L2[4][23+1], L1[13][23], L1[13+1][23], L1[13+2][23]);

assign L2[5][24] = L1[0][24];
fa fa_L2_66(L2[6][24], L2[0][24+1], L1[1][24], L1[1+1][24], L1[1+2][24]);
fa fa_L2_67(L2[7][24], L2[1][24+1], L1[4][24], L1[4+1][24], L1[4+2][24]);
fa fa_L2_68(L2[8][24], L2[2][24+1], L1[7][24], L1[7+1][24], L1[7+2][24]);
fa fa_L2_69(L2[9][24], L2[3][24+1], L1[10][24], L1[10+1][24], L1[10+2][24]);
fa fa_L2_70(L2[10][24], L2[4][24+1], L1[13][24], L1[13+1][24], L1[13+2][24]);

assign L2[5][25] = L1[0][25];
fa fa_L2_71(L2[6][25], L2[0][25+1], L1[1][25], L1[1+1][25], L1[1+2][25]);
fa fa_L2_72(L2[7][25], L2[1][25+1], L1[4][25], L1[4+1][25], L1[4+2][25]);
fa fa_L2_73(L2[8][25], L2[2][25+1], L1[7][25], L1[7+1][25], L1[7+2][25]);
fa fa_L2_74(L2[9][25], L2[3][25+1], L1[10][25], L1[10+1][25], L1[10+2][25]);
fa fa_L2_75(L2[10][25], L2[4][25+1], L1[13][25], L1[13+1][25], L1[13+2][25]);

ha ha_L2_76(L2[5][26], L2[0][26+1], L1[0][26], L1[0+1][26]);
fa fa_L2_77(L2[6][26], L2[1][26+1], L1[2][26], L1[2+1][26], L1[2+2][26]);
fa fa_L2_78(L2[7][26], L2[2][26+1], L1[5][26], L1[5+1][26], L1[5+2][26]);
fa fa_L2_79(L2[8][26], L2[3][26+1], L1[8][26], L1[8+1][26], L1[8+2][26]);
fa fa_L2_80(L2[9][26], L2[4][26+1], L1[11][26], L1[11+1][26], L1[11+2][26]);

ha ha_L2_81(L2[5][27], L2[0][27+1], L1[0][27], L1[0+1][27]);
fa fa_L2_82(L2[6][27], L2[1][27+1], L1[2][27], L1[2+1][27], L1[2+2][27]);
fa fa_L2_83(L2[7][27], L2[2][27+1], L1[5][27], L1[5+1][27], L1[5+2][27]);
fa fa_L2_84(L2[8][27], L2[3][27+1], L1[8][27], L1[8+1][27], L1[8+2][27]);
fa fa_L2_85(L2[9][27], L2[4][27+1], L1[11][27], L1[11+1][27], L1[11+2][27]);

ha ha_L2_86(L2[5][28], L2[0][28+1], L1[0][28], L1[0+1][28]);
fa fa_L2_87(L2[6][28], L2[1][28+1], L1[2][28], L1[2+1][28], L1[2+2][28]);
fa fa_L2_88(L2[7][28], L2[2][28+1], L1[5][28], L1[5+1][28], L1[5+2][28]);
fa fa_L2_89(L2[8][28], L2[3][28+1], L1[8][28], L1[8+1][28], L1[8+2][28]);
fa fa_L2_90(L2[9][28], L2[4][28+1], L1[11][28], L1[11+1][28], L1[11+2][28]);

fa fa_L2_91(L2[5][29], L2[0][29+1], L1[0][29], L1[0+1][29], L1[0+2][29]);
fa fa_L2_92(L2[6][29], L2[1][29+1], L1[3][29], L1[3+1][29], L1[3+2][29]);
fa fa_L2_93(L2[7][29], L2[2][29+1], L1[6][29], L1[6+1][29], L1[6+2][29]);
fa fa_L2_94(L2[8][29], L2[3][29+1], L1[9][29], L1[9+1][29], L1[9+2][29]);

fa fa_L2_95(L2[4][30], L2[0][30+1], L1[0][30], L1[0+1][30], L1[0+2][30]);
fa fa_L2_96(L2[5][30], L2[1][30+1], L1[3][30], L1[3+1][30], L1[3+2][30]);
fa fa_L2_97(L2[6][30], L2[2][30+1], L1[6][30], L1[6+1][30], L1[6+2][30]);
fa fa_L2_98(L2[7][30], L2[3][30+1], L1[9][30], L1[9+1][30], L1[9+2][30]);

fa fa_L2_99(L2[4][31], L2[0][31+1], L1[0][31], L1[0+1][31], L1[0+2][31]);
fa fa_L2_100(L2[5][31], L2[1][31+1], L1[3][31], L1[3+1][31], L1[3+2][31]);
fa fa_L2_101(L2[6][31], L2[2][31+1], L1[6][31], L1[6+1][31], L1[6+2][31]);
fa fa_L2_102(L2[7][31], L2[3][31+1], L1[9][31], L1[9+1][31], L1[9+2][31]);

assign L2[4][32] = L1[0][32];
fa fa_L2_103(L2[5][32], L2[0][32+1], L1[1][32], L1[1+1][32], L1[1+2][32]);
fa fa_L2_104(L2[6][32], L2[1][32+1], L1[4][32], L1[4+1][32], L1[4+2][32]);
fa fa_L2_105(L2[7][32], L2[2][32+1], L1[7][32], L1[7+1][32], L1[7+2][32]);

assign L2[3][33] = L1[0][33];
fa fa_L2_106(L2[4][33], L2[0][33+1], L1[1][33], L1[1+1][33], L1[1+2][33]);
fa fa_L2_107(L2[5][33], L2[1][33+1], L1[4][33], L1[4+1][33], L1[4+2][33]);
fa fa_L2_108(L2[6][33], L2[2][33+1], L1[7][33], L1[7+1][33], L1[7+2][33]);

assign L2[3][34] = L1[0][34];
fa fa_L2_109(L2[4][34], L2[0][34+1], L1[1][34], L1[1+1][34], L1[1+2][34]);
fa fa_L2_110(L2[5][34], L2[1][34+1], L1[4][34], L1[4+1][34], L1[4+2][34]);
fa fa_L2_111(L2[6][34], L2[2][34+1], L1[7][34], L1[7+1][34], L1[7+2][34]);

ha ha_L2_112(L2[3][35], L2[0][35+1], L1[0][35], L1[0+1][35]);
fa fa_L2_113(L2[4][35], L2[1][35+1], L1[2][35], L1[2+1][35], L1[2+2][35]);
fa fa_L2_114(L2[5][35], L2[2][35+1], L1[5][35], L1[5+1][35], L1[5+2][35]);

ha ha_L2_115(L2[3][36], L2[0][36+1], L1[0][36], L1[0+1][36]);
fa fa_L2_116(L2[4][36], L2[1][36+1], L1[2][36], L1[2+1][36], L1[2+2][36]);
fa fa_L2_117(L2[5][36], L2[2][36+1], L1[5][36], L1[5+1][36], L1[5+2][36]);

ha ha_L2_118(L2[3][37], L2[0][37+1], L1[0][37], L1[0+1][37]);
fa fa_L2_119(L2[4][37], L2[1][37+1], L1[2][37], L1[2+1][37], L1[2+2][37]);
fa fa_L2_120(L2[5][37], L2[2][37+1], L1[5][37], L1[5+1][37], L1[5+2][37]);

fa fa_L2_121(L2[3][38], L2[0][38+1], L1[0][38], L1[0+1][38], L1[0+2][38]);
fa fa_L2_122(L2[4][38], L2[1][38+1], L1[3][38], L1[3+1][38], L1[3+2][38]);

fa fa_L2_123(L2[2][39], L2[0][39+1], L1[0][39], L1[0+1][39], L1[0+2][39]);
fa fa_L2_124(L2[3][39], L2[1][39+1], L1[3][39], L1[3+1][39], L1[3+2][39]);

fa fa_L2_125(L2[2][40], L2[0][40+1], L1[0][40], L1[0+1][40], L1[0+2][40]);
fa fa_L2_126(L2[3][40], L2[1][40+1], L1[3][40], L1[3+1][40], L1[3+2][40]);

assign L2[2][41] = L1[0][41];
fa fa_L2_127(L2[3][41], L2[0][41+1], L1[1][41], L1[1+1][41], L1[1+2][41]);

assign L2[1][42] = L1[0][42];
fa fa_L2_128(L2[2][42], L2[0][42+1], L1[1][42], L1[1+1][42], L1[1+2][42]);

assign L2[1][43] = L1[0][43];
fa fa_L2_129(L2[2][43], L2[0][43+1], L1[1][43], L1[1+1][43], L1[1+2][43]);

ha ha_L2_130(L2[1][44], L2[0][44+1], L1[0][44], L1[0+1][44]);

fa fa_L2_131(L2[1][45], L2[0][45+1], L1[0][45], L1[0+1][45], L1[0+2][45]);

assign L2[1][46] = L1[0][46];


assign L3[0][0] = L2[0][0];

assign L3[0][1] = L2[0][1];

assign L3[0][2] = L2[0][2];

ha ha_L3_0(L3[0][3], L3[0][3+1], L2[0][3], L2[0+1][3]);

ha ha_L3_1(L3[1][4], L3[0][4+1], L2[0][4], L2[0+1][4]);

fa fa_L3_2(L3[1][5], L3[0][5+1], L2[0][5], L2[0+1][5], L2[0+2][5]);

fa fa_L3_3(L3[1][6], L3[0][6+1], L2[0][6], L2[0+1][6], L2[0+2][6]);

assign L3[1][7] = L2[0][7];
fa fa_L3_4(L3[2][7], L3[0][7+1], L2[1][7], L2[1+1][7], L2[1+2][7]);

assign L3[1][8] = L2[0][8];
fa fa_L3_5(L3[2][8], L3[0][8+1], L2[1][8], L2[1+1][8], L2[1+2][8]);

ha ha_L3_6(L3[1][9], L3[0][9+1], L2[0][9], L2[0+1][9]);
fa fa_L3_7(L3[2][9], L3[1][9+1], L2[2][9], L2[2+1][9], L2[2+2][9]);

ha ha_L3_8(L3[2][10], L3[0][10+1], L2[0][10], L2[0+1][10]);
fa fa_L3_9(L3[3][10], L3[1][10+1], L2[2][10], L2[2+1][10], L2[2+2][10]);

ha ha_L3_10(L3[2][11], L3[0][11+1], L2[0][11], L2[0+1][11]);
fa fa_L3_11(L3[3][11], L3[1][11+1], L2[2][11], L2[2+1][11], L2[2+2][11]);

fa fa_L3_12(L3[2][12], L3[0][12+1], L2[0][12], L2[0+1][12], L2[0+2][12]);
fa fa_L3_13(L3[3][12], L3[1][12+1], L2[3][12], L2[3+1][12], L2[3+2][12]);

fa fa_L3_14(L3[2][13], L3[0][13+1], L2[0][13], L2[0+1][13], L2[0+2][13]);
fa fa_L3_15(L3[3][13], L3[1][13+1], L2[3][13], L2[3+1][13], L2[3+2][13]);

assign L3[2][14] = L2[0][14];
fa fa_L3_16(L3[3][14], L3[0][14+1], L2[1][14], L2[1+1][14], L2[1+2][14]);
fa fa_L3_17(L3[4][14], L3[1][14+1], L2[4][14], L2[4+1][14], L2[4+2][14]);

assign L3[2][15] = L2[0][15];
fa fa_L3_18(L3[3][15], L3[0][15+1], L2[1][15], L2[1+1][15], L2[1+2][15]);
fa fa_L3_19(L3[4][15], L3[1][15+1], L2[4][15], L2[4+1][15], L2[4+2][15]);

ha ha_L3_20(L3[2][16], L3[0][16+1], L2[0][16], L2[0+1][16]);
fa fa_L3_21(L3[3][16], L3[1][16+1], L2[2][16], L2[2+1][16], L2[2+2][16]);
fa fa_L3_22(L3[4][16], L3[2][16+1], L2[5][16], L2[5+1][16], L2[5+2][16]);

ha ha_L3_23(L3[3][17], L3[0][17+1], L2[0][17], L2[0+1][17]);
fa fa_L3_24(L3[4][17], L3[1][17+1], L2[2][17], L2[2+1][17], L2[2+2][17]);
fa fa_L3_25(L3[5][17], L3[2][17+1], L2[5][17], L2[5+1][17], L2[5+2][17]);

fa fa_L3_26(L3[3][18], L3[0][18+1], L2[0][18], L2[0+1][18], L2[0+2][18]);
fa fa_L3_27(L3[4][18], L3[1][18+1], L2[3][18], L2[3+1][18], L2[3+2][18]);
fa fa_L3_28(L3[5][18], L3[2][18+1], L2[6][18], L2[6+1][18], L2[6+2][18]);

fa fa_L3_29(L3[3][19], L3[0][19+1], L2[0][19], L2[0+1][19], L2[0+2][19]);
fa fa_L3_30(L3[4][19], L3[1][19+1], L2[3][19], L2[3+1][19], L2[3+2][19]);
fa fa_L3_31(L3[5][19], L3[2][19+1], L2[6][19], L2[6+1][19], L2[6+2][19]);

fa fa_L3_32(L3[3][20], L3[0][20+1], L2[0][20], L2[0+1][20], L2[0+2][20]);
fa fa_L3_33(L3[4][20], L3[1][20+1], L2[3][20], L2[3+1][20], L2[3+2][20]);
fa fa_L3_34(L3[5][20], L3[2][20+1], L2[6][20], L2[6+1][20], L2[6+2][20]);

assign L3[3][21] = L2[0][21];
fa fa_L3_35(L3[4][21], L3[0][21+1], L2[1][21], L2[1+1][21], L2[1+2][21]);
fa fa_L3_36(L3[5][21], L3[1][21+1], L2[4][21], L2[4+1][21], L2[4+2][21]);
fa fa_L3_37(L3[6][21], L3[2][21+1], L2[7][21], L2[7+1][21], L2[7+2][21]);

assign L3[3][22] = L2[0][22];
fa fa_L3_38(L3[4][22], L3[0][22+1], L2[1][22], L2[1+1][22], L2[1+2][22]);
fa fa_L3_39(L3[5][22], L3[1][22+1], L2[4][22], L2[4+1][22], L2[4+2][22]);
fa fa_L3_40(L3[6][22], L3[2][22+1], L2[7][22], L2[7+1][22], L2[7+2][22]);

ha ha_L3_41(L3[3][23], L3[0][23+1], L2[0][23], L2[0+1][23]);
fa fa_L3_42(L3[4][23], L3[1][23+1], L2[2][23], L2[2+1][23], L2[2+2][23]);
fa fa_L3_43(L3[5][23], L3[2][23+1], L2[5][23], L2[5+1][23], L2[5+2][23]);
fa fa_L3_44(L3[6][23], L3[3][23+1], L2[8][23], L2[8+1][23], L2[8+2][23]);

ha ha_L3_45(L3[4][24], L3[0][24+1], L2[0][24], L2[0+1][24]);
fa fa_L3_46(L3[5][24], L3[1][24+1], L2[2][24], L2[2+1][24], L2[2+2][24]);
fa fa_L3_47(L3[6][24], L3[2][24+1], L2[5][24], L2[5+1][24], L2[5+2][24]);
fa fa_L3_48(L3[7][24], L3[3][24+1], L2[8][24], L2[8+1][24], L2[8+2][24]);

ha ha_L3_49(L3[4][25], L3[0][25+1], L2[0][25], L2[0+1][25]);
fa fa_L3_50(L3[5][25], L3[1][25+1], L2[2][25], L2[2+1][25], L2[2+2][25]);
fa fa_L3_51(L3[6][25], L3[2][25+1], L2[5][25], L2[5+1][25], L2[5+2][25]);
fa fa_L3_52(L3[7][25], L3[3][25+1], L2[8][25], L2[8+1][25], L2[8+2][25]);

assign L3[4][26] = L2[0][26];
fa fa_L3_53(L3[5][26], L3[0][26+1], L2[1][26], L2[1+1][26], L2[1+2][26]);
fa fa_L3_54(L3[6][26], L3[1][26+1], L2[4][26], L2[4+1][26], L2[4+2][26]);
fa fa_L3_55(L3[7][26], L3[2][26+1], L2[7][26], L2[7+1][26], L2[7+2][26]);

assign L3[3][27] = L2[0][27];
fa fa_L3_56(L3[4][27], L3[0][27+1], L2[1][27], L2[1+1][27], L2[1+2][27]);
fa fa_L3_57(L3[5][27], L3[1][27+1], L2[4][27], L2[4+1][27], L2[4+2][27]);
fa fa_L3_58(L3[6][27], L3[2][27+1], L2[7][27], L2[7+1][27], L2[7+2][27]);

assign L3[3][28] = L2[0][28];
fa fa_L3_59(L3[4][28], L3[0][28+1], L2[1][28], L2[1+1][28], L2[1+2][28]);
fa fa_L3_60(L3[5][28], L3[1][28+1], L2[4][28], L2[4+1][28], L2[4+2][28]);
fa fa_L3_61(L3[6][28], L3[2][28+1], L2[7][28], L2[7+1][28], L2[7+2][28]);

fa fa_L3_62(L3[3][29], L3[0][29+1], L2[0][29], L2[0+1][29], L2[0+2][29]);
fa fa_L3_63(L3[4][29], L3[1][29+1], L2[3][29], L2[3+1][29], L2[3+2][29]);
fa fa_L3_64(L3[5][29], L3[2][29+1], L2[6][29], L2[6+1][29], L2[6+2][29]);

ha ha_L3_65(L3[3][30], L3[0][30+1], L2[0][30], L2[0+1][30]);
fa fa_L3_66(L3[4][30], L3[1][30+1], L2[2][30], L2[2+1][30], L2[2+2][30]);
fa fa_L3_67(L3[5][30], L3[2][30+1], L2[5][30], L2[5+1][30], L2[5+2][30]);

ha ha_L3_68(L3[3][31], L3[0][31+1], L2[0][31], L2[0+1][31]);
fa fa_L3_69(L3[4][31], L3[1][31+1], L2[2][31], L2[2+1][31], L2[2+2][31]);
fa fa_L3_70(L3[5][31], L3[2][31+1], L2[5][31], L2[5+1][31], L2[5+2][31]);

ha ha_L3_71(L3[3][32], L3[0][32+1], L2[0][32], L2[0+1][32]);
fa fa_L3_72(L3[4][32], L3[1][32+1], L2[2][32], L2[2+1][32], L2[2+2][32]);
fa fa_L3_73(L3[5][32], L3[2][32+1], L2[5][32], L2[5+1][32], L2[5+2][32]);

assign L3[3][33] = L2[0][33];
fa fa_L3_74(L3[4][33], L3[0][33+1], L2[1][33], L2[1+1][33], L2[1+2][33]);
fa fa_L3_75(L3[5][33], L3[1][33+1], L2[4][33], L2[4+1][33], L2[4+2][33]);

assign L3[2][34] = L2[0][34];
fa fa_L3_76(L3[3][34], L3[0][34+1], L2[1][34], L2[1+1][34], L2[1+2][34]);
fa fa_L3_77(L3[4][34], L3[1][34+1], L2[4][34], L2[4+1][34], L2[4+2][34]);

fa fa_L3_78(L3[2][35], L3[0][35+1], L2[0][35], L2[0+1][35], L2[0+2][35]);
fa fa_L3_79(L3[3][35], L3[1][35+1], L2[3][35], L2[3+1][35], L2[3+2][35]);

fa fa_L3_80(L3[2][36], L3[0][36+1], L2[0][36], L2[0+1][36], L2[0+2][36]);
fa fa_L3_81(L3[3][36], L3[1][36+1], L2[3][36], L2[3+1][36], L2[3+2][36]);

fa fa_L3_82(L3[2][37], L3[0][37+1], L2[0][37], L2[0+1][37], L2[0+2][37]);
fa fa_L3_83(L3[3][37], L3[1][37+1], L2[3][37], L2[3+1][37], L2[3+2][37]);

ha ha_L3_84(L3[2][38], L3[0][38+1], L2[0][38], L2[0+1][38]);
fa fa_L3_85(L3[3][38], L3[1][38+1], L2[2][38], L2[2+1][38], L2[2+2][38]);

assign L3[2][39] = L2[0][39];
fa fa_L3_86(L3[3][39], L3[0][39+1], L2[1][39], L2[1+1][39], L2[1+2][39]);

assign L3[1][40] = L2[0][40];
fa fa_L3_87(L3[2][40], L3[0][40+1], L2[1][40], L2[1+1][40], L2[1+2][40]);

assign L3[1][41] = L2[0][41];
fa fa_L3_88(L3[2][41], L3[0][41+1], L2[1][41], L2[1+1][41], L2[1+2][41]);

fa fa_L3_89(L3[1][42], L3[0][42+1], L2[0][42], L2[0+1][42], L2[0+2][42]);

fa fa_L3_90(L3[1][43], L3[0][43+1], L2[0][43], L2[0+1][43], L2[0+2][43]);

assign L3[1][44] = L2[0][44];
assign L3[2][44] = L2[1][44];

assign L3[0][45] = L2[0][45];
assign L3[1][45] = L2[1][45];

assign L3[0][46] = L2[0][46];
assign L3[1][46] = L2[1][46];


assign L4[0][0] = L3[0][0];

assign L4[0][1] = L3[0][1];

assign L4[0][2] = L3[0][2];

assign L4[0][3] = L3[0][3];

ha ha_L4_0(L4[0][4], L4[0][4+1], L3[0][4], L3[0+1][4]);

ha ha_L4_1(L4[1][5], L4[0][5+1], L3[0][5], L3[0+1][5]);

ha ha_L4_2(L4[1][6], L4[0][6+1], L3[0][6], L3[0+1][6]);

fa fa_L4_3(L4[1][7], L4[0][7+1], L3[0][7], L3[0+1][7], L3[0+2][7]);

fa fa_L4_4(L4[1][8], L4[0][8+1], L3[0][8], L3[0+1][8], L3[0+2][8]);

fa fa_L4_5(L4[1][9], L4[0][9+1], L3[0][9], L3[0+1][9], L3[0+2][9]);

assign L4[1][10] = L3[0][10];
fa fa_L4_6(L4[2][10], L4[0][10+1], L3[1][10], L3[1+1][10], L3[1+2][10]);

assign L4[1][11] = L3[0][11];
fa fa_L4_7(L4[2][11], L4[0][11+1], L3[1][11], L3[1+1][11], L3[1+2][11]);

assign L4[1][12] = L3[0][12];
fa fa_L4_8(L4[2][12], L4[0][12+1], L3[1][12], L3[1+1][12], L3[1+2][12]);

assign L4[1][13] = L3[0][13];
fa fa_L4_9(L4[2][13], L4[0][13+1], L3[1][13], L3[1+1][13], L3[1+2][13]);

ha ha_L4_10(L4[1][14], L4[0][14+1], L3[0][14], L3[0+1][14]);
fa fa_L4_11(L4[2][14], L4[1][14+1], L3[2][14], L3[2+1][14], L3[2+2][14]);

ha ha_L4_12(L4[2][15], L4[0][15+1], L3[0][15], L3[0+1][15]);
fa fa_L4_13(L4[3][15], L4[1][15+1], L3[2][15], L3[2+1][15], L3[2+2][15]);

ha ha_L4_14(L4[2][16], L4[0][16+1], L3[0][16], L3[0+1][16]);
fa fa_L4_15(L4[3][16], L4[1][16+1], L3[2][16], L3[2+1][16], L3[2+2][16]);

fa fa_L4_16(L4[2][17], L4[0][17+1], L3[0][17], L3[0+1][17], L3[0+2][17]);
fa fa_L4_17(L4[3][17], L4[1][17+1], L3[3][17], L3[3+1][17], L3[3+2][17]);

fa fa_L4_18(L4[2][18], L4[0][18+1], L3[0][18], L3[0+1][18], L3[0+2][18]);
fa fa_L4_19(L4[3][18], L4[1][18+1], L3[3][18], L3[3+1][18], L3[3+2][18]);

fa fa_L4_20(L4[2][19], L4[0][19+1], L3[0][19], L3[0+1][19], L3[0+2][19]);
fa fa_L4_21(L4[3][19], L4[1][19+1], L3[3][19], L3[3+1][19], L3[3+2][19]);

fa fa_L4_22(L4[2][20], L4[0][20+1], L3[0][20], L3[0+1][20], L3[0+2][20]);
fa fa_L4_23(L4[3][20], L4[1][20+1], L3[3][20], L3[3+1][20], L3[3+2][20]);

assign L4[2][21] = L3[0][21];
fa fa_L4_24(L4[3][21], L4[0][21+1], L3[1][21], L3[1+1][21], L3[1+2][21]);
fa fa_L4_25(L4[4][21], L4[1][21+1], L3[4][21], L3[4+1][21], L3[4+2][21]);

assign L4[2][22] = L3[0][22];
fa fa_L4_26(L4[3][22], L4[0][22+1], L3[1][22], L3[1+1][22], L3[1+2][22]);
fa fa_L4_27(L4[4][22], L4[1][22+1], L3[4][22], L3[4+1][22], L3[4+2][22]);

assign L4[2][23] = L3[0][23];
fa fa_L4_28(L4[3][23], L4[0][23+1], L3[1][23], L3[1+1][23], L3[1+2][23]);
fa fa_L4_29(L4[4][23], L4[1][23+1], L3[4][23], L3[4+1][23], L3[4+2][23]);

ha ha_L4_30(L4[2][24], L4[0][24+1], L3[0][24], L3[0+1][24]);
fa fa_L4_31(L4[3][24], L4[1][24+1], L3[2][24], L3[2+1][24], L3[2+2][24]);
fa fa_L4_32(L4[4][24], L4[2][24+1], L3[5][24], L3[5+1][24], L3[5+2][24]);

ha ha_L4_33(L4[3][25], L4[0][25+1], L3[0][25], L3[0+1][25]);
fa fa_L4_34(L4[4][25], L4[1][25+1], L3[2][25], L3[2+1][25], L3[2+2][25]);
fa fa_L4_35(L4[5][25], L4[2][25+1], L3[5][25], L3[5+1][25], L3[5+2][25]);

ha ha_L4_36(L4[3][26], L4[0][26+1], L3[0][26], L3[0+1][26]);
fa fa_L4_37(L4[4][26], L4[1][26+1], L3[2][26], L3[2+1][26], L3[2+2][26]);
fa fa_L4_38(L4[5][26], L4[2][26+1], L3[5][26], L3[5+1][26], L3[5+2][26]);

assign L4[3][27] = L3[0][27];
fa fa_L4_39(L4[4][27], L4[0][27+1], L3[1][27], L3[1+1][27], L3[1+2][27]);
fa fa_L4_40(L4[5][27], L4[1][27+1], L3[4][27], L3[4+1][27], L3[4+2][27]);

assign L4[2][28] = L3[0][28];
fa fa_L4_41(L4[3][28], L4[0][28+1], L3[1][28], L3[1+1][28], L3[1+2][28]);
fa fa_L4_42(L4[4][28], L4[1][28+1], L3[4][28], L3[4+1][28], L3[4+2][28]);

fa fa_L4_43(L4[2][29], L4[0][29+1], L3[0][29], L3[0+1][29], L3[0+2][29]);
fa fa_L4_44(L4[3][29], L4[1][29+1], L3[3][29], L3[3+1][29], L3[3+2][29]);

fa fa_L4_45(L4[2][30], L4[0][30+1], L3[0][30], L3[0+1][30], L3[0+2][30]);
fa fa_L4_46(L4[3][30], L4[1][30+1], L3[3][30], L3[3+1][30], L3[3+2][30]);

fa fa_L4_47(L4[2][31], L4[0][31+1], L3[0][31], L3[0+1][31], L3[0+2][31]);
fa fa_L4_48(L4[3][31], L4[1][31+1], L3[3][31], L3[3+1][31], L3[3+2][31]);

fa fa_L4_49(L4[2][32], L4[0][32+1], L3[0][32], L3[0+1][32], L3[0+2][32]);
fa fa_L4_50(L4[3][32], L4[1][32+1], L3[3][32], L3[3+1][32], L3[3+2][32]);

fa fa_L4_51(L4[2][33], L4[0][33+1], L3[0][33], L3[0+1][33], L3[0+2][33]);
fa fa_L4_52(L4[3][33], L4[1][33+1], L3[3][33], L3[3+1][33], L3[3+2][33]);

ha ha_L4_53(L4[2][34], L4[0][34+1], L3[0][34], L3[0+1][34]);
fa fa_L4_54(L4[3][34], L4[1][34+1], L3[2][34], L3[2+1][34], L3[2+2][34]);

assign L4[2][35] = L3[0][35];
fa fa_L4_55(L4[3][35], L4[0][35+1], L3[1][35], L3[1+1][35], L3[1+2][35]);

assign L4[1][36] = L3[0][36];
fa fa_L4_56(L4[2][36], L4[0][36+1], L3[1][36], L3[1+1][36], L3[1+2][36]);

assign L4[1][37] = L3[0][37];
fa fa_L4_57(L4[2][37], L4[0][37+1], L3[1][37], L3[1+1][37], L3[1+2][37]);

assign L4[1][38] = L3[0][38];
fa fa_L4_58(L4[2][38], L4[0][38+1], L3[1][38], L3[1+1][38], L3[1+2][38]);

assign L4[1][39] = L3[0][39];
fa fa_L4_59(L4[2][39], L4[0][39+1], L3[1][39], L3[1+1][39], L3[1+2][39]);

fa fa_L4_60(L4[1][40], L4[0][40+1], L3[0][40], L3[0+1][40], L3[0+2][40]);

fa fa_L4_61(L4[1][41], L4[0][41+1], L3[0][41], L3[0+1][41], L3[0+2][41]);

ha ha_L4_62(L4[1][42], L4[0][42+1], L3[0][42], L3[0+1][42]);

ha ha_L4_63(L4[1][43], L4[0][43+1], L3[0][43], L3[0+1][43]);

fa fa_L4_64(L4[1][44], L4[0][44+1], L3[0][44], L3[0+1][44], L3[0+2][44]);

assign L4[1][45] = L3[0][45];
assign L4[2][45] = L3[1][45];

assign L4[0][46] = L3[0][46];
assign L4[1][46] = L3[1][46];


assign L5[0][0] = L4[0][0];

assign L5[0][1] = L4[0][1];

assign L5[0][2] = L4[0][2];

assign L5[0][3] = L4[0][3];

assign L5[0][4] = L4[0][4];

ha ha_L5_0(L5[0][5], L5[0][5+1], L4[0][5], L4[0+1][5]);

ha ha_L5_1(L5[1][6], L5[0][6+1], L4[0][6], L4[0+1][6]);

ha ha_L5_2(L5[1][7], L5[0][7+1], L4[0][7], L4[0+1][7]);

ha ha_L5_3(L5[1][8], L5[0][8+1], L4[0][8], L4[0+1][8]);

ha ha_L5_4(L5[1][9], L5[0][9+1], L4[0][9], L4[0+1][9]);

fa fa_L5_5(L5[1][10], L5[0][10+1], L4[0][10], L4[0+1][10], L4[0+2][10]);

fa fa_L5_6(L5[1][11], L5[0][11+1], L4[0][11], L4[0+1][11], L4[0+2][11]);

fa fa_L5_7(L5[1][12], L5[0][12+1], L4[0][12], L4[0+1][12], L4[0+2][12]);

fa fa_L5_8(L5[1][13], L5[0][13+1], L4[0][13], L4[0+1][13], L4[0+2][13]);

fa fa_L5_9(L5[1][14], L5[0][14+1], L4[0][14], L4[0+1][14], L4[0+2][14]);

assign L5[1][15] = L4[0][15];
fa fa_L5_10(L5[2][15], L5[0][15+1], L4[1][15], L4[1+1][15], L4[1+2][15]);

assign L5[1][16] = L4[0][16];
fa fa_L5_11(L5[2][16], L5[0][16+1], L4[1][16], L4[1+1][16], L4[1+2][16]);

assign L5[1][17] = L4[0][17];
fa fa_L5_12(L5[2][17], L5[0][17+1], L4[1][17], L4[1+1][17], L4[1+2][17]);

assign L5[1][18] = L4[0][18];
fa fa_L5_13(L5[2][18], L5[0][18+1], L4[1][18], L4[1+1][18], L4[1+2][18]);

assign L5[1][19] = L4[0][19];
fa fa_L5_14(L5[2][19], L5[0][19+1], L4[1][19], L4[1+1][19], L4[1+2][19]);

assign L5[1][20] = L4[0][20];
fa fa_L5_15(L5[2][20], L5[0][20+1], L4[1][20], L4[1+1][20], L4[1+2][20]);

ha ha_L5_16(L5[1][21], L5[0][21+1], L4[0][21], L4[0+1][21]);
fa fa_L5_17(L5[2][21], L5[1][21+1], L4[2][21], L4[2+1][21], L4[2+2][21]);

ha ha_L5_18(L5[2][22], L5[0][22+1], L4[0][22], L4[0+1][22]);
fa fa_L5_19(L5[3][22], L5[1][22+1], L4[2][22], L4[2+1][22], L4[2+2][22]);

ha ha_L5_20(L5[2][23], L5[0][23+1], L4[0][23], L4[0+1][23]);
fa fa_L5_21(L5[3][23], L5[1][23+1], L4[2][23], L4[2+1][23], L4[2+2][23]);

ha ha_L5_22(L5[2][24], L5[0][24+1], L4[0][24], L4[0+1][24]);
fa fa_L5_23(L5[3][24], L5[1][24+1], L4[2][24], L4[2+1][24], L4[2+2][24]);

fa fa_L5_24(L5[2][25], L5[0][25+1], L4[0][25], L4[0+1][25], L4[0+2][25]);
fa fa_L5_25(L5[3][25], L5[1][25+1], L4[3][25], L4[3+1][25], L4[3+2][25]);

fa fa_L5_26(L5[2][26], L5[0][26+1], L4[0][26], L4[0+1][26], L4[0+2][26]);
fa fa_L5_27(L5[3][26], L5[1][26+1], L4[3][26], L4[3+1][26], L4[3+2][26]);

fa fa_L5_28(L5[2][27], L5[0][27+1], L4[0][27], L4[0+1][27], L4[0+2][27]);
fa fa_L5_29(L5[3][27], L5[1][27+1], L4[3][27], L4[3+1][27], L4[3+2][27]);

ha ha_L5_30(L5[2][28], L5[0][28+1], L4[0][28], L4[0+1][28]);
fa fa_L5_31(L5[3][28], L5[1][28+1], L4[2][28], L4[2+1][28], L4[2+2][28]);

assign L5[2][29] = L4[0][29];
fa fa_L5_32(L5[3][29], L5[0][29+1], L4[1][29], L4[1+1][29], L4[1+2][29]);

assign L5[1][30] = L4[0][30];
fa fa_L5_33(L5[2][30], L5[0][30+1], L4[1][30], L4[1+1][30], L4[1+2][30]);

assign L5[1][31] = L4[0][31];
fa fa_L5_34(L5[2][31], L5[0][31+1], L4[1][31], L4[1+1][31], L4[1+2][31]);

assign L5[1][32] = L4[0][32];
fa fa_L5_35(L5[2][32], L5[0][32+1], L4[1][32], L4[1+1][32], L4[1+2][32]);

assign L5[1][33] = L4[0][33];
fa fa_L5_36(L5[2][33], L5[0][33+1], L4[1][33], L4[1+1][33], L4[1+2][33]);

assign L5[1][34] = L4[0][34];
fa fa_L5_37(L5[2][34], L5[0][34+1], L4[1][34], L4[1+1][34], L4[1+2][34]);

assign L5[1][35] = L4[0][35];
fa fa_L5_38(L5[2][35], L5[0][35+1], L4[1][35], L4[1+1][35], L4[1+2][35]);

fa fa_L5_39(L5[1][36], L5[0][36+1], L4[0][36], L4[0+1][36], L4[0+2][36]);

fa fa_L5_40(L5[1][37], L5[0][37+1], L4[0][37], L4[0+1][37], L4[0+2][37]);

fa fa_L5_41(L5[1][38], L5[0][38+1], L4[0][38], L4[0+1][38], L4[0+2][38]);

fa fa_L5_42(L5[1][39], L5[0][39+1], L4[0][39], L4[0+1][39], L4[0+2][39]);

ha ha_L5_43(L5[1][40], L5[0][40+1], L4[0][40], L4[0+1][40]);

ha ha_L5_44(L5[1][41], L5[0][41+1], L4[0][41], L4[0+1][41]);

ha ha_L5_45(L5[1][42], L5[0][42+1], L4[0][42], L4[0+1][42]);

ha ha_L5_46(L5[1][43], L5[0][43+1], L4[0][43], L4[0+1][43]);

ha ha_L5_47(L5[1][44], L5[0][44+1], L4[0][44], L4[0+1][44]);

fa fa_L5_48(L5[1][45], L5[0][45+1], L4[0][45], L4[0+1][45], L4[0+2][45]);

assign L5[1][46] = L4[0][46];
assign L5[2][46] = L4[1][46];


assign L6[0][0] = L5[0][0];

assign L6[0][1] = L5[0][1];

assign L6[0][2] = L5[0][2];

assign L6[0][3] = L5[0][3];

assign L6[0][4] = L5[0][4];

assign L6[0][5] = L5[0][5];

ha ha_L6_0(L6[0][6], L6[0][6+1], L5[0][6], L5[0+1][6]);

ha ha_L6_1(L6[1][7], L6[0][7+1], L5[0][7], L5[0+1][7]);

ha ha_L6_2(L6[1][8], L6[0][8+1], L5[0][8], L5[0+1][8]);

ha ha_L6_3(L6[1][9], L6[0][9+1], L5[0][9], L5[0+1][9]);

ha ha_L6_4(L6[1][10], L6[0][10+1], L5[0][10], L5[0+1][10]);

ha ha_L6_5(L6[1][11], L6[0][11+1], L5[0][11], L5[0+1][11]);

ha ha_L6_6(L6[1][12], L6[0][12+1], L5[0][12], L5[0+1][12]);

ha ha_L6_7(L6[1][13], L6[0][13+1], L5[0][13], L5[0+1][13]);

ha ha_L6_8(L6[1][14], L6[0][14+1], L5[0][14], L5[0+1][14]);

fa fa_L6_9(L6[1][15], L6[0][15+1], L5[0][15], L5[0+1][15], L5[0+2][15]);

fa fa_L6_10(L6[1][16], L6[0][16+1], L5[0][16], L5[0+1][16], L5[0+2][16]);

fa fa_L6_11(L6[1][17], L6[0][17+1], L5[0][17], L5[0+1][17], L5[0+2][17]);

fa fa_L6_12(L6[1][18], L6[0][18+1], L5[0][18], L5[0+1][18], L5[0+2][18]);

fa fa_L6_13(L6[1][19], L6[0][19+1], L5[0][19], L5[0+1][19], L5[0+2][19]);

fa fa_L6_14(L6[1][20], L6[0][20+1], L5[0][20], L5[0+1][20], L5[0+2][20]);

fa fa_L6_15(L6[1][21], L6[0][21+1], L5[0][21], L5[0+1][21], L5[0+2][21]);

assign L6[1][22] = L5[0][22];
fa fa_L6_16(L6[2][22], L6[0][22+1], L5[1][22], L5[1+1][22], L5[1+2][22]);

assign L6[1][23] = L5[0][23];
fa fa_L6_17(L6[2][23], L6[0][23+1], L5[1][23], L5[1+1][23], L5[1+2][23]);

assign L6[1][24] = L5[0][24];
fa fa_L6_18(L6[2][24], L6[0][24+1], L5[1][24], L5[1+1][24], L5[1+2][24]);

assign L6[1][25] = L5[0][25];
fa fa_L6_19(L6[2][25], L6[0][25+1], L5[1][25], L5[1+1][25], L5[1+2][25]);

assign L6[1][26] = L5[0][26];
fa fa_L6_20(L6[2][26], L6[0][26+1], L5[1][26], L5[1+1][26], L5[1+2][26]);

assign L6[1][27] = L5[0][27];
fa fa_L6_21(L6[2][27], L6[0][27+1], L5[1][27], L5[1+1][27], L5[1+2][27]);

assign L6[1][28] = L5[0][28];
fa fa_L6_22(L6[2][28], L6[0][28+1], L5[1][28], L5[1+1][28], L5[1+2][28]);

assign L6[1][29] = L5[0][29];
fa fa_L6_23(L6[2][29], L6[0][29+1], L5[1][29], L5[1+1][29], L5[1+2][29]);

fa fa_L6_24(L6[1][30], L6[0][30+1], L5[0][30], L5[0+1][30], L5[0+2][30]);

fa fa_L6_25(L6[1][31], L6[0][31+1], L5[0][31], L5[0+1][31], L5[0+2][31]);

fa fa_L6_26(L6[1][32], L6[0][32+1], L5[0][32], L5[0+1][32], L5[0+2][32]);

fa fa_L6_27(L6[1][33], L6[0][33+1], L5[0][33], L5[0+1][33], L5[0+2][33]);

fa fa_L6_28(L6[1][34], L6[0][34+1], L5[0][34], L5[0+1][34], L5[0+2][34]);

fa fa_L6_29(L6[1][35], L6[0][35+1], L5[0][35], L5[0+1][35], L5[0+2][35]);

ha ha_L6_30(L6[1][36], L6[0][36+1], L5[0][36], L5[0+1][36]);

ha ha_L6_31(L6[1][37], L6[0][37+1], L5[0][37], L5[0+1][37]);

ha ha_L6_32(L6[1][38], L6[0][38+1], L5[0][38], L5[0+1][38]);

ha ha_L6_33(L6[1][39], L6[0][39+1], L5[0][39], L5[0+1][39]);

ha ha_L6_34(L6[1][40], L6[0][40+1], L5[0][40], L5[0+1][40]);

ha ha_L6_35(L6[1][41], L6[0][41+1], L5[0][41], L5[0+1][41]);

ha ha_L6_36(L6[1][42], L6[0][42+1], L5[0][42], L5[0+1][42]);

ha ha_L6_37(L6[1][43], L6[0][43+1], L5[0][43], L5[0+1][43]);

ha ha_L6_38(L6[1][44], L6[0][44+1], L5[0][44], L5[0+1][44]);

ha ha_L6_39(L6[1][45], L6[0][45+1], L5[0][45], L5[0+1][45]);

fa fa_L6_40(L6[1][46], L6[0][46+1], L5[0][46], L5[0+1][46], L5[0+2][46]);


assign L7[0][0] = L6[0][0];

assign L7[0][1] = L6[0][1];

assign L7[0][2] = L6[0][2];

assign L7[0][3] = L6[0][3];

assign L7[0][4] = L6[0][4];

assign L7[0][5] = L6[0][5];

assign L7[0][6] = L6[0][6];

ha ha_L7_0(L7[0][7], L7[0][7+1], L6[0][7], L6[0+1][7]);

ha ha_L7_1(L7[1][8], L7[0][8+1], L6[0][8], L6[0+1][8]);

ha ha_L7_2(L7[1][9], L7[0][9+1], L6[0][9], L6[0+1][9]);

ha ha_L7_3(L7[1][10], L7[0][10+1], L6[0][10], L6[0+1][10]);

ha ha_L7_4(L7[1][11], L7[0][11+1], L6[0][11], L6[0+1][11]);

ha ha_L7_5(L7[1][12], L7[0][12+1], L6[0][12], L6[0+1][12]);

ha ha_L7_6(L7[1][13], L7[0][13+1], L6[0][13], L6[0+1][13]);

ha ha_L7_7(L7[1][14], L7[0][14+1], L6[0][14], L6[0+1][14]);

ha ha_L7_8(L7[1][15], L7[0][15+1], L6[0][15], L6[0+1][15]);

ha ha_L7_9(L7[1][16], L7[0][16+1], L6[0][16], L6[0+1][16]);

ha ha_L7_10(L7[1][17], L7[0][17+1], L6[0][17], L6[0+1][17]);

ha ha_L7_11(L7[1][18], L7[0][18+1], L6[0][18], L6[0+1][18]);

ha ha_L7_12(L7[1][19], L7[0][19+1], L6[0][19], L6[0+1][19]);

ha ha_L7_13(L7[1][20], L7[0][20+1], L6[0][20], L6[0+1][20]);

ha ha_L7_14(L7[1][21], L7[0][21+1], L6[0][21], L6[0+1][21]);

fa fa_L7_15(L7[1][22], L7[0][22+1], L6[0][22], L6[0+1][22], L6[0+2][22]);

fa fa_L7_16(L7[1][23], L7[0][23+1], L6[0][23], L6[0+1][23], L6[0+2][23]);

fa fa_L7_17(L7[1][24], L7[0][24+1], L6[0][24], L6[0+1][24], L6[0+2][24]);

fa fa_L7_18(L7[1][25], L7[0][25+1], L6[0][25], L6[0+1][25], L6[0+2][25]);

fa fa_L7_19(L7[1][26], L7[0][26+1], L6[0][26], L6[0+1][26], L6[0+2][26]);

fa fa_L7_20(L7[1][27], L7[0][27+1], L6[0][27], L6[0+1][27], L6[0+2][27]);

fa fa_L7_21(L7[1][28], L7[0][28+1], L6[0][28], L6[0+1][28], L6[0+2][28]);

fa fa_L7_22(L7[1][29], L7[0][29+1], L6[0][29], L6[0+1][29], L6[0+2][29]);

ha ha_L7_23(L7[1][30], L7[0][30+1], L6[0][30], L6[0+1][30]);

ha ha_L7_24(L7[1][31], L7[0][31+1], L6[0][31], L6[0+1][31]);

ha ha_L7_25(L7[1][32], L7[0][32+1], L6[0][32], L6[0+1][32]);

ha ha_L7_26(L7[1][33], L7[0][33+1], L6[0][33], L6[0+1][33]);

ha ha_L7_27(L7[1][34], L7[0][34+1], L6[0][34], L6[0+1][34]);

ha ha_L7_28(L7[1][35], L7[0][35+1], L6[0][35], L6[0+1][35]);

ha ha_L7_29(L7[1][36], L7[0][36+1], L6[0][36], L6[0+1][36]);

ha ha_L7_30(L7[1][37], L7[0][37+1], L6[0][37], L6[0+1][37]);

ha ha_L7_31(L7[1][38], L7[0][38+1], L6[0][38], L6[0+1][38]);

ha ha_L7_32(L7[1][39], L7[0][39+1], L6[0][39], L6[0+1][39]);

ha ha_L7_33(L7[1][40], L7[0][40+1], L6[0][40], L6[0+1][40]);

ha ha_L7_34(L7[1][41], L7[0][41+1], L6[0][41], L6[0+1][41]);

ha ha_L7_35(L7[1][42], L7[0][42+1], L6[0][42], L6[0+1][42]);

ha ha_L7_36(L7[1][43], L7[0][43+1], L6[0][43], L6[0+1][43]);

ha ha_L7_37(L7[1][44], L7[0][44+1], L6[0][44], L6[0+1][44]);

ha ha_L7_38(L7[1][45], L7[0][45+1], L6[0][45], L6[0+1][45]);

ha ha_L7_39(L7[1][46], L7[0][46+1], L6[0][46], L6[0+1][46]);

assign L7[1][47] = L6[0][47];



endmodule
