// Dadda mult
module dadda_mult(
    output [47:0] product,
    input [23:0] A, B
);

wire [46:0] partial_products[23:0];

// i=1, j=23 => 1-(1+23-23)
// Partial product generation
genvar i, j;
generate
    for (i = 0; i < 24; i = i + 1) begin : pp_generation
        for (j = 0; j < 24; j = j + 1) begin : pp_gen
            if(i+j>23) begin  //If column idx is larger than bit width,
                assign partial_products[23-j][i+j] = A[j] & B[i];
            end
            else begin
                assign partial_products[i][i+j] = A[j] & B[i];
            end
        end
    end
endgenerate

wire [47:0] L1[22:0];
wire [47:0] L2[22:0];
wire [47:0] L3[22:0];
wire [47:0] L4[22:0];
wire [47:0] L5[22:0];
wire [47:0] L6[22:0];
wire [47:0] L7[22:0];

//45-bit adder
assign product[0] = L7[0][0];
adder adder_inst(
    .A(L7[0][46:1]),
    .B(L7[1][46:1]), 
    .Sum(product[46:1]), 
    .Cout(product[47])
    );

assign L1[0][0] = partial_products[0][0];

assign L1[0][1] = partial_products[0][1];
assign L1[1][1] = partial_products[1][1];

assign L1[0][2] = partial_products[0][2];
assign L1[1][2] = partial_products[1][2];
assign L1[2][2] = partial_products[2][2];

assign L1[0][3] = partial_products[0][3];
assign L1[1][3] = partial_products[1][3];
assign L1[2][3] = partial_products[2][3];
assign L1[3][3] = partial_products[3][3];

assign L1[0][4] = partial_products[0][4];
assign L1[1][4] = partial_products[1][4];
assign L1[2][4] = partial_products[2][4];
assign L1[3][4] = partial_products[3][4];
assign L1[4][4] = partial_products[4][4];

assign L1[0][5] = partial_products[0][5];
assign L1[1][5] = partial_products[1][5];
assign L1[2][5] = partial_products[2][5];
assign L1[3][5] = partial_products[3][5];
assign L1[4][5] = partial_products[4][5];
assign L1[5][5] = partial_products[5][5];

assign L1[0][6] = partial_products[0][6];
assign L1[1][6] = partial_products[1][6];
assign L1[2][6] = partial_products[2][6];
assign L1[3][6] = partial_products[3][6];
assign L1[4][6] = partial_products[4][6];
assign L1[5][6] = partial_products[5][6];
assign L1[6][6] = partial_products[6][6];

assign L1[0][7] = partial_products[0][7];
assign L1[1][7] = partial_products[1][7];
assign L1[2][7] = partial_products[2][7];
assign L1[3][7] = partial_products[3][7];
assign L1[4][7] = partial_products[4][7];
assign L1[5][7] = partial_products[5][7];
assign L1[6][7] = partial_products[6][7];
assign L1[7][7] = partial_products[7][7];

assign L1[0][8] = partial_products[0][8];
assign L1[1][8] = partial_products[1][8];
assign L1[2][8] = partial_products[2][8];
assign L1[3][8] = partial_products[3][8];
assign L1[4][8] = partial_products[4][8];
assign L1[5][8] = partial_products[5][8];
assign L1[6][8] = partial_products[6][8];
assign L1[7][8] = partial_products[7][8];
assign L1[8][8] = partial_products[8][8];

assign L1[0][9] = partial_products[0][9];
assign L1[1][9] = partial_products[1][9];
assign L1[2][9] = partial_products[2][9];
assign L1[3][9] = partial_products[3][9];
assign L1[4][9] = partial_products[4][9];
assign L1[5][9] = partial_products[5][9];
assign L1[6][9] = partial_products[6][9];
assign L1[7][9] = partial_products[7][9];
assign L1[8][9] = partial_products[8][9];
assign L1[9][9] = partial_products[9][9];

assign L1[0][10] = partial_products[0][10];
assign L1[1][10] = partial_products[1][10];
assign L1[2][10] = partial_products[2][10];
assign L1[3][10] = partial_products[3][10];
assign L1[4][10] = partial_products[4][10];
assign L1[5][10] = partial_products[5][10];
assign L1[6][10] = partial_products[6][10];
assign L1[7][10] = partial_products[7][10];
assign L1[8][10] = partial_products[8][10];
assign L1[9][10] = partial_products[9][10];
assign L1[10][10] = partial_products[10][10];

assign L1[0][11] = partial_products[0][11];
assign L1[1][11] = partial_products[1][11];
assign L1[2][11] = partial_products[2][11];
assign L1[3][11] = partial_products[3][11];
assign L1[4][11] = partial_products[4][11];
assign L1[5][11] = partial_products[5][11];
assign L1[6][11] = partial_products[6][11];
assign L1[7][11] = partial_products[7][11];
assign L1[8][11] = partial_products[8][11];
assign L1[9][11] = partial_products[9][11];
assign L1[10][11] = partial_products[10][11];
assign L1[11][11] = partial_products[11][11];

assign L1[0][12] = partial_products[0][12];
assign L1[1][12] = partial_products[1][12];
assign L1[2][12] = partial_products[2][12];
assign L1[3][12] = partial_products[3][12];
assign L1[4][12] = partial_products[4][12];
assign L1[5][12] = partial_products[5][12];
assign L1[6][12] = partial_products[6][12];
assign L1[7][12] = partial_products[7][12];
assign L1[8][12] = partial_products[8][12];
assign L1[9][12] = partial_products[9][12];
assign L1[10][12] = partial_products[10][12];
assign L1[11][12] = partial_products[11][12];
assign L1[12][12] = partial_products[12][12];

assign L1[0][13] = partial_products[0][13];
assign L1[1][13] = partial_products[1][13];
assign L1[2][13] = partial_products[2][13];
assign L1[3][13] = partial_products[3][13];
assign L1[4][13] = partial_products[4][13];
assign L1[5][13] = partial_products[5][13];
assign L1[6][13] = partial_products[6][13];
assign L1[7][13] = partial_products[7][13];
assign L1[8][13] = partial_products[8][13];
assign L1[9][13] = partial_products[9][13];
assign L1[10][13] = partial_products[10][13];
assign L1[11][13] = partial_products[11][13];
assign L1[12][13] = partial_products[12][13];
assign L1[13][13] = partial_products[13][13];

assign L1[0][14] = partial_products[0][14];
assign L1[1][14] = partial_products[1][14];
assign L1[2][14] = partial_products[2][14];
assign L1[3][14] = partial_products[3][14];
assign L1[4][14] = partial_products[4][14];
assign L1[5][14] = partial_products[5][14];
assign L1[6][14] = partial_products[6][14];
assign L1[7][14] = partial_products[7][14];
assign L1[8][14] = partial_products[8][14];
assign L1[9][14] = partial_products[9][14];
assign L1[10][14] = partial_products[10][14];
assign L1[11][14] = partial_products[11][14];
assign L1[12][14] = partial_products[12][14];
assign L1[13][14] = partial_products[13][14];
assign L1[14][14] = partial_products[14][14];

assign L1[0][15] = partial_products[0][15];
assign L1[1][15] = partial_products[1][15];
assign L1[2][15] = partial_products[2][15];
assign L1[3][15] = partial_products[3][15];
assign L1[4][15] = partial_products[4][15];
assign L1[5][15] = partial_products[5][15];
assign L1[6][15] = partial_products[6][15];
assign L1[7][15] = partial_products[7][15];
assign L1[8][15] = partial_products[8][15];
assign L1[9][15] = partial_products[9][15];
assign L1[10][15] = partial_products[10][15];
assign L1[11][15] = partial_products[11][15];
assign L1[12][15] = partial_products[12][15];
assign L1[13][15] = partial_products[13][15];
assign L1[14][15] = partial_products[14][15];
assign L1[15][15] = partial_products[15][15];

assign L1[0][16] = partial_products[0][16];
assign L1[1][16] = partial_products[1][16];
assign L1[2][16] = partial_products[2][16];
assign L1[3][16] = partial_products[3][16];
assign L1[4][16] = partial_products[4][16];
assign L1[5][16] = partial_products[5][16];
assign L1[6][16] = partial_products[6][16];
assign L1[7][16] = partial_products[7][16];
assign L1[8][16] = partial_products[8][16];
assign L1[9][16] = partial_products[9][16];
assign L1[10][16] = partial_products[10][16];
assign L1[11][16] = partial_products[11][16];
assign L1[12][16] = partial_products[12][16];
assign L1[13][16] = partial_products[13][16];
assign L1[14][16] = partial_products[14][16];
assign L1[15][16] = partial_products[15][16];
assign L1[16][16] = partial_products[16][16];

assign L1[0][17] = partial_products[0][17];
assign L1[1][17] = partial_products[1][17];
assign L1[2][17] = partial_products[2][17];
assign L1[3][17] = partial_products[3][17];
assign L1[4][17] = partial_products[4][17];
assign L1[5][17] = partial_products[5][17];
assign L1[6][17] = partial_products[6][17];
assign L1[7][17] = partial_products[7][17];
assign L1[8][17] = partial_products[8][17];
assign L1[9][17] = partial_products[9][17];
assign L1[10][17] = partial_products[10][17];
assign L1[11][17] = partial_products[11][17];
assign L1[12][17] = partial_products[12][17];
assign L1[13][17] = partial_products[13][17];
assign L1[14][17] = partial_products[14][17];
assign L1[15][17] = partial_products[15][17];
assign L1[16][17] = partial_products[16][17];
assign L1[17][17] = partial_products[17][17];

assign L1[0][18] = partial_products[0][18];
assign L1[1][18] = partial_products[1][18];
assign L1[2][18] = partial_products[2][18];
assign L1[3][18] = partial_products[3][18];
assign L1[4][18] = partial_products[4][18];
assign L1[5][18] = partial_products[5][18];
assign L1[6][18] = partial_products[6][18];
assign L1[7][18] = partial_products[7][18];
assign L1[8][18] = partial_products[8][18];
assign L1[9][18] = partial_products[9][18];
assign L1[10][18] = partial_products[10][18];
assign L1[11][18] = partial_products[11][18];
assign L1[12][18] = partial_products[12][18];
assign L1[13][18] = partial_products[13][18];
assign L1[14][18] = partial_products[14][18];
assign L1[15][18] = partial_products[15][18];
assign L1[16][18] = partial_products[16][18];
assign L1[17][18] = partial_products[17][18];
assign L1[18][18] = partial_products[18][18];

assign { L1[0][19+1], L1[0][19] } = partial_products[0][19] + partial_products[0+1][19];
assign L1[1][19] = partial_products[2][19];
assign L1[2][19] = partial_products[3][19];
assign L1[3][19] = partial_products[4][19];
assign L1[4][19] = partial_products[5][19];
assign L1[5][19] = partial_products[6][19];
assign L1[6][19] = partial_products[7][19];
assign L1[7][19] = partial_products[8][19];
assign L1[8][19] = partial_products[9][19];
assign L1[9][19] = partial_products[10][19];
assign L1[10][19] = partial_products[11][19];
assign L1[11][19] = partial_products[12][19];
assign L1[12][19] = partial_products[13][19];
assign L1[13][19] = partial_products[14][19];
assign L1[14][19] = partial_products[15][19];
assign L1[15][19] = partial_products[16][19];
assign L1[16][19] = partial_products[17][19];
assign L1[17][19] = partial_products[18][19];
assign L1[18][19] = partial_products[19][19];

assign { L1[0][20+1], L1[1][20] } = partial_products[0][20] + partial_products[0+1][20] + partial_products[0+2][20];
assign { L1[1][20+1], L1[2][20] } = partial_products[3][20] + partial_products[3+1][20];
assign L1[3][20] = partial_products[5][20];
assign L1[4][20] = partial_products[6][20];
assign L1[5][20] = partial_products[7][20];
assign L1[6][20] = partial_products[8][20];
assign L1[7][20] = partial_products[9][20];
assign L1[8][20] = partial_products[10][20];
assign L1[9][20] = partial_products[11][20];
assign L1[10][20] = partial_products[12][20];
assign L1[11][20] = partial_products[13][20];
assign L1[12][20] = partial_products[14][20];
assign L1[13][20] = partial_products[15][20];
assign L1[14][20] = partial_products[16][20];
assign L1[15][20] = partial_products[17][20];
assign L1[16][20] = partial_products[18][20];
assign L1[17][20] = partial_products[19][20];
assign L1[18][20] = partial_products[20][20];

assign { L1[0][21+1], L1[2][21] } = partial_products[0][21] + partial_products[0+1][21] + partial_products[0+2][21];
assign { L1[1][21+1], L1[3][21] } = partial_products[3][21] + partial_products[3+1][21] + partial_products[3+2][21];
assign { L1[2][21+1], L1[4][21] } = partial_products[6][21] + partial_products[6+1][21];
assign L1[5][21] = partial_products[8][21];
assign L1[6][21] = partial_products[9][21];
assign L1[7][21] = partial_products[10][21];
assign L1[8][21] = partial_products[11][21];
assign L1[9][21] = partial_products[12][21];
assign L1[10][21] = partial_products[13][21];
assign L1[11][21] = partial_products[14][21];
assign L1[12][21] = partial_products[15][21];
assign L1[13][21] = partial_products[16][21];
assign L1[14][21] = partial_products[17][21];
assign L1[15][21] = partial_products[18][21];
assign L1[16][21] = partial_products[19][21];
assign L1[17][21] = partial_products[20][21];
assign L1[18][21] = partial_products[21][21];

assign { L1[0][22+1], L1[3][22] } = partial_products[0][22] + partial_products[0+1][22] + partial_products[0+2][22];
assign { L1[1][22+1], L1[4][22] } = partial_products[3][22] + partial_products[3+1][22] + partial_products[3+2][22];
assign { L1[2][22+1], L1[5][22] } = partial_products[6][22] + partial_products[6+1][22] + partial_products[6+2][22];
assign { L1[3][22+1], L1[6][22] } = partial_products[9][22] + partial_products[9+1][22];
assign L1[7][22] = partial_products[11][22];
assign L1[8][22] = partial_products[12][22];
assign L1[9][22] = partial_products[13][22];
assign L1[10][22] = partial_products[14][22];
assign L1[11][22] = partial_products[15][22];
assign L1[12][22] = partial_products[16][22];
assign L1[13][22] = partial_products[17][22];
assign L1[14][22] = partial_products[18][22];
assign L1[15][22] = partial_products[19][22];
assign L1[16][22] = partial_products[20][22];
assign L1[17][22] = partial_products[21][22];
assign L1[18][22] = partial_products[22][22];

assign { L1[0][23+1], L1[4][23] } = partial_products[0][23] + partial_products[0+1][23] + partial_products[0+2][23];
assign { L1[1][23+1], L1[5][23] } = partial_products[3][23] + partial_products[3+1][23] + partial_products[3+2][23];
assign { L1[2][23+1], L1[6][23] } = partial_products[6][23] + partial_products[6+1][23] + partial_products[6+2][23];
assign { L1[3][23+1], L1[7][23] } = partial_products[9][23] + partial_products[9+1][23] + partial_products[9+2][23];
assign { L1[4][23+1], L1[8][23] } = partial_products[12][23] + partial_products[12+1][23];
assign L1[9][23] = partial_products[14][23];
assign L1[10][23] = partial_products[15][23];
assign L1[11][23] = partial_products[16][23];
assign L1[12][23] = partial_products[17][23];
assign L1[13][23] = partial_products[18][23];
assign L1[14][23] = partial_products[19][23];
assign L1[15][23] = partial_products[20][23];
assign L1[16][23] = partial_products[21][23];
assign L1[17][23] = partial_products[22][23];
assign L1[18][23] = partial_products[23][23];

assign { L1[0][24+1], L1[5][24] } = partial_products[0][24] + partial_products[0+1][24] + partial_products[0+2][24];
assign { L1[1][24+1], L1[6][24] } = partial_products[3][24] + partial_products[3+1][24] + partial_products[3+2][24];
assign { L1[2][24+1], L1[7][24] } = partial_products[6][24] + partial_products[6+1][24] + partial_products[6+2][24];
assign { L1[3][24+1], L1[8][24] } = partial_products[9][24] + partial_products[9+1][24] + partial_products[9+2][24];
assign { L1[4][24+1], L1[9][24] } = partial_products[12][24] + partial_products[12+1][24];
assign L1[10][24] = partial_products[14][24];
assign L1[11][24] = partial_products[15][24];
assign L1[12][24] = partial_products[16][24];
assign L1[13][24] = partial_products[17][24];
assign L1[14][24] = partial_products[18][24];
assign L1[15][24] = partial_products[19][24];
assign L1[16][24] = partial_products[20][24];
assign L1[17][24] = partial_products[21][24];
assign L1[18][24] = partial_products[22][24];

assign { L1[0][25+1], L1[5][25] } = partial_products[0][25] + partial_products[0+1][25] + partial_products[0+2][25];
assign { L1[1][25+1], L1[6][25] } = partial_products[3][25] + partial_products[3+1][25] + partial_products[3+2][25];
assign { L1[2][25+1], L1[7][25] } = partial_products[6][25] + partial_products[6+1][25] + partial_products[6+2][25];
assign { L1[3][25+1], L1[8][25] } = partial_products[9][25] + partial_products[9+1][25] + partial_products[9+2][25];
assign L1[9][25] = partial_products[12][25];
assign L1[10][25] = partial_products[13][25];
assign L1[11][25] = partial_products[14][25];
assign L1[12][25] = partial_products[15][25];
assign L1[13][25] = partial_products[16][25];
assign L1[14][25] = partial_products[17][25];
assign L1[15][25] = partial_products[18][25];
assign L1[16][25] = partial_products[19][25];
assign L1[17][25] = partial_products[20][25];
assign L1[18][25] = partial_products[21][25];

assign { L1[0][26+1], L1[4][26] } = partial_products[0][26] + partial_products[0+1][26] + partial_products[0+2][26];
assign { L1[1][26+1], L1[5][26] } = partial_products[3][26] + partial_products[3+1][26] + partial_products[3+2][26];
assign { L1[2][26+1], L1[6][26] } = partial_products[6][26] + partial_products[6+1][26] + partial_products[6+2][26];
assign L1[7][26] = partial_products[9][26];
assign L1[8][26] = partial_products[10][26];
assign L1[9][26] = partial_products[11][26];
assign L1[10][26] = partial_products[12][26];
assign L1[11][26] = partial_products[13][26];
assign L1[12][26] = partial_products[14][26];
assign L1[13][26] = partial_products[15][26];
assign L1[14][26] = partial_products[16][26];
assign L1[15][26] = partial_products[17][26];
assign L1[16][26] = partial_products[18][26];
assign L1[17][26] = partial_products[19][26];
assign L1[18][26] = partial_products[20][26];

assign { L1[0][27+1], L1[3][27] } = partial_products[0][27] + partial_products[0+1][27] + partial_products[0+2][27];
assign { L1[1][27+1], L1[4][27] } = partial_products[3][27] + partial_products[3+1][27] + partial_products[3+2][27];
assign L1[5][27] = partial_products[6][27];
assign L1[6][27] = partial_products[7][27];
assign L1[7][27] = partial_products[8][27];
assign L1[8][27] = partial_products[9][27];
assign L1[9][27] = partial_products[10][27];
assign L1[10][27] = partial_products[11][27];
assign L1[11][27] = partial_products[12][27];
assign L1[12][27] = partial_products[13][27];
assign L1[13][27] = partial_products[14][27];
assign L1[14][27] = partial_products[15][27];
assign L1[15][27] = partial_products[16][27];
assign L1[16][27] = partial_products[17][27];
assign L1[17][27] = partial_products[18][27];
assign L1[18][27] = partial_products[19][27];

assign { L1[0][28+1], L1[2][28] } = partial_products[0][28] + partial_products[0+1][28] + partial_products[0+2][28];
assign L1[3][28] = partial_products[3][28];
assign L1[4][28] = partial_products[4][28];
assign L1[5][28] = partial_products[5][28];
assign L1[6][28] = partial_products[6][28];
assign L1[7][28] = partial_products[7][28];
assign L1[8][28] = partial_products[8][28];
assign L1[9][28] = partial_products[9][28];
assign L1[10][28] = partial_products[10][28];
assign L1[11][28] = partial_products[11][28];
assign L1[12][28] = partial_products[12][28];
assign L1[13][28] = partial_products[13][28];
assign L1[14][28] = partial_products[14][28];
assign L1[15][28] = partial_products[15][28];
assign L1[16][28] = partial_products[16][28];
assign L1[17][28] = partial_products[17][28];
assign L1[18][28] = partial_products[18][28];

assign L1[1][29] = partial_products[0][29];
assign L1[2][29] = partial_products[1][29];
assign L1[3][29] = partial_products[2][29];
assign L1[4][29] = partial_products[3][29];
assign L1[5][29] = partial_products[4][29];
assign L1[6][29] = partial_products[5][29];
assign L1[7][29] = partial_products[6][29];
assign L1[8][29] = partial_products[7][29];
assign L1[9][29] = partial_products[8][29];
assign L1[10][29] = partial_products[9][29];
assign L1[11][29] = partial_products[10][29];
assign L1[12][29] = partial_products[11][29];
assign L1[13][29] = partial_products[12][29];
assign L1[14][29] = partial_products[13][29];
assign L1[15][29] = partial_products[14][29];
assign L1[16][29] = partial_products[15][29];
assign L1[17][29] = partial_products[16][29];
assign L1[18][29] = partial_products[17][29];

assign L1[0][30] = partial_products[0][30];
assign L1[1][30] = partial_products[1][30];
assign L1[2][30] = partial_products[2][30];
assign L1[3][30] = partial_products[3][30];
assign L1[4][30] = partial_products[4][30];
assign L1[5][30] = partial_products[5][30];
assign L1[6][30] = partial_products[6][30];
assign L1[7][30] = partial_products[7][30];
assign L1[8][30] = partial_products[8][30];
assign L1[9][30] = partial_products[9][30];
assign L1[10][30] = partial_products[10][30];
assign L1[11][30] = partial_products[11][30];
assign L1[12][30] = partial_products[12][30];
assign L1[13][30] = partial_products[13][30];
assign L1[14][30] = partial_products[14][30];
assign L1[15][30] = partial_products[15][30];
assign L1[16][30] = partial_products[16][30];

assign L1[0][31] = partial_products[0][31];
assign L1[1][31] = partial_products[1][31];
assign L1[2][31] = partial_products[2][31];
assign L1[3][31] = partial_products[3][31];
assign L1[4][31] = partial_products[4][31];
assign L1[5][31] = partial_products[5][31];
assign L1[6][31] = partial_products[6][31];
assign L1[7][31] = partial_products[7][31];
assign L1[8][31] = partial_products[8][31];
assign L1[9][31] = partial_products[9][31];
assign L1[10][31] = partial_products[10][31];
assign L1[11][31] = partial_products[11][31];
assign L1[12][31] = partial_products[12][31];
assign L1[13][31] = partial_products[13][31];
assign L1[14][31] = partial_products[14][31];
assign L1[15][31] = partial_products[15][31];

assign L1[0][32] = partial_products[0][32];
assign L1[1][32] = partial_products[1][32];
assign L1[2][32] = partial_products[2][32];
assign L1[3][32] = partial_products[3][32];
assign L1[4][32] = partial_products[4][32];
assign L1[5][32] = partial_products[5][32];
assign L1[6][32] = partial_products[6][32];
assign L1[7][32] = partial_products[7][32];
assign L1[8][32] = partial_products[8][32];
assign L1[9][32] = partial_products[9][32];
assign L1[10][32] = partial_products[10][32];
assign L1[11][32] = partial_products[11][32];
assign L1[12][32] = partial_products[12][32];
assign L1[13][32] = partial_products[13][32];
assign L1[14][32] = partial_products[14][32];

assign L1[0][33] = partial_products[0][33];
assign L1[1][33] = partial_products[1][33];
assign L1[2][33] = partial_products[2][33];
assign L1[3][33] = partial_products[3][33];
assign L1[4][33] = partial_products[4][33];
assign L1[5][33] = partial_products[5][33];
assign L1[6][33] = partial_products[6][33];
assign L1[7][33] = partial_products[7][33];
assign L1[8][33] = partial_products[8][33];
assign L1[9][33] = partial_products[9][33];
assign L1[10][33] = partial_products[10][33];
assign L1[11][33] = partial_products[11][33];
assign L1[12][33] = partial_products[12][33];
assign L1[13][33] = partial_products[13][33];

assign L1[0][34] = partial_products[0][34];
assign L1[1][34] = partial_products[1][34];
assign L1[2][34] = partial_products[2][34];
assign L1[3][34] = partial_products[3][34];
assign L1[4][34] = partial_products[4][34];
assign L1[5][34] = partial_products[5][34];
assign L1[6][34] = partial_products[6][34];
assign L1[7][34] = partial_products[7][34];
assign L1[8][34] = partial_products[8][34];
assign L1[9][34] = partial_products[9][34];
assign L1[10][34] = partial_products[10][34];
assign L1[11][34] = partial_products[11][34];
assign L1[12][34] = partial_products[12][34];

assign L1[0][35] = partial_products[0][35];
assign L1[1][35] = partial_products[1][35];
assign L1[2][35] = partial_products[2][35];
assign L1[3][35] = partial_products[3][35];
assign L1[4][35] = partial_products[4][35];
assign L1[5][35] = partial_products[5][35];
assign L1[6][35] = partial_products[6][35];
assign L1[7][35] = partial_products[7][35];
assign L1[8][35] = partial_products[8][35];
assign L1[9][35] = partial_products[9][35];
assign L1[10][35] = partial_products[10][35];
assign L1[11][35] = partial_products[11][35];

assign L1[0][36] = partial_products[0][36];
assign L1[1][36] = partial_products[1][36];
assign L1[2][36] = partial_products[2][36];
assign L1[3][36] = partial_products[3][36];
assign L1[4][36] = partial_products[4][36];
assign L1[5][36] = partial_products[5][36];
assign L1[6][36] = partial_products[6][36];
assign L1[7][36] = partial_products[7][36];
assign L1[8][36] = partial_products[8][36];
assign L1[9][36] = partial_products[9][36];
assign L1[10][36] = partial_products[10][36];

assign L1[0][37] = partial_products[0][37];
assign L1[1][37] = partial_products[1][37];
assign L1[2][37] = partial_products[2][37];
assign L1[3][37] = partial_products[3][37];
assign L1[4][37] = partial_products[4][37];
assign L1[5][37] = partial_products[5][37];
assign L1[6][37] = partial_products[6][37];
assign L1[7][37] = partial_products[7][37];
assign L1[8][37] = partial_products[8][37];
assign L1[9][37] = partial_products[9][37];

assign L1[0][38] = partial_products[0][38];
assign L1[1][38] = partial_products[1][38];
assign L1[2][38] = partial_products[2][38];
assign L1[3][38] = partial_products[3][38];
assign L1[4][38] = partial_products[4][38];
assign L1[5][38] = partial_products[5][38];
assign L1[6][38] = partial_products[6][38];
assign L1[7][38] = partial_products[7][38];
assign L1[8][38] = partial_products[8][38];

assign L1[0][39] = partial_products[0][39];
assign L1[1][39] = partial_products[1][39];
assign L1[2][39] = partial_products[2][39];
assign L1[3][39] = partial_products[3][39];
assign L1[4][39] = partial_products[4][39];
assign L1[5][39] = partial_products[5][39];
assign L1[6][39] = partial_products[6][39];
assign L1[7][39] = partial_products[7][39];

assign L1[0][40] = partial_products[0][40];
assign L1[1][40] = partial_products[1][40];
assign L1[2][40] = partial_products[2][40];
assign L1[3][40] = partial_products[3][40];
assign L1[4][40] = partial_products[4][40];
assign L1[5][40] = partial_products[5][40];
assign L1[6][40] = partial_products[6][40];

assign L1[0][41] = partial_products[0][41];
assign L1[1][41] = partial_products[1][41];
assign L1[2][41] = partial_products[2][41];
assign L1[3][41] = partial_products[3][41];
assign L1[4][41] = partial_products[4][41];
assign L1[5][41] = partial_products[5][41];

assign L1[0][42] = partial_products[0][42];
assign L1[1][42] = partial_products[1][42];
assign L1[2][42] = partial_products[2][42];
assign L1[3][42] = partial_products[3][42];
assign L1[4][42] = partial_products[4][42];

assign L1[0][43] = partial_products[0][43];
assign L1[1][43] = partial_products[1][43];
assign L1[2][43] = partial_products[2][43];
assign L1[3][43] = partial_products[3][43];

assign L1[0][44] = partial_products[0][44];
assign L1[1][44] = partial_products[1][44];
assign L1[2][44] = partial_products[2][44];

assign L1[0][45] = partial_products[0][45];
assign L1[1][45] = partial_products[1][45];

assign L1[0][46] = partial_products[0][46];


assign L2[0][0] = L1[0][0];

assign L2[0][1] = L1[0][1];
assign L2[1][1] = L1[1][1];

assign L2[0][2] = L1[0][2];
assign L2[1][2] = L1[1][2];
assign L2[2][2] = L1[2][2];

assign L2[0][3] = L1[0][3];
assign L2[1][3] = L1[1][3];
assign L2[2][3] = L1[2][3];
assign L2[3][3] = L1[3][3];

assign L2[0][4] = L1[0][4];
assign L2[1][4] = L1[1][4];
assign L2[2][4] = L1[2][4];
assign L2[3][4] = L1[3][4];
assign L2[4][4] = L1[4][4];

assign L2[0][5] = L1[0][5];
assign L2[1][5] = L1[1][5];
assign L2[2][5] = L1[2][5];
assign L2[3][5] = L1[3][5];
assign L2[4][5] = L1[4][5];
assign L2[5][5] = L1[5][5];

assign L2[0][6] = L1[0][6];
assign L2[1][6] = L1[1][6];
assign L2[2][6] = L1[2][6];
assign L2[3][6] = L1[3][6];
assign L2[4][6] = L1[4][6];
assign L2[5][6] = L1[5][6];
assign L2[6][6] = L1[6][6];

assign L2[0][7] = L1[0][7];
assign L2[1][7] = L1[1][7];
assign L2[2][7] = L1[2][7];
assign L2[3][7] = L1[3][7];
assign L2[4][7] = L1[4][7];
assign L2[5][7] = L1[5][7];
assign L2[6][7] = L1[6][7];
assign L2[7][7] = L1[7][7];

assign L2[0][8] = L1[0][8];
assign L2[1][8] = L1[1][8];
assign L2[2][8] = L1[2][8];
assign L2[3][8] = L1[3][8];
assign L2[4][8] = L1[4][8];
assign L2[5][8] = L1[5][8];
assign L2[6][8] = L1[6][8];
assign L2[7][8] = L1[7][8];
assign L2[8][8] = L1[8][8];

assign L2[0][9] = L1[0][9];
assign L2[1][9] = L1[1][9];
assign L2[2][9] = L1[2][9];
assign L2[3][9] = L1[3][9];
assign L2[4][9] = L1[4][9];
assign L2[5][9] = L1[5][9];
assign L2[6][9] = L1[6][9];
assign L2[7][9] = L1[7][9];
assign L2[8][9] = L1[8][9];
assign L2[9][9] = L1[9][9];

assign L2[0][10] = L1[0][10];
assign L2[1][10] = L1[1][10];
assign L2[2][10] = L1[2][10];
assign L2[3][10] = L1[3][10];
assign L2[4][10] = L1[4][10];
assign L2[5][10] = L1[5][10];
assign L2[6][10] = L1[6][10];
assign L2[7][10] = L1[7][10];
assign L2[8][10] = L1[8][10];
assign L2[9][10] = L1[9][10];
assign L2[10][10] = L1[10][10];

assign L2[0][11] = L1[0][11];
assign L2[1][11] = L1[1][11];
assign L2[2][11] = L1[2][11];
assign L2[3][11] = L1[3][11];
assign L2[4][11] = L1[4][11];
assign L2[5][11] = L1[5][11];
assign L2[6][11] = L1[6][11];
assign L2[7][11] = L1[7][11];
assign L2[8][11] = L1[8][11];
assign L2[9][11] = L1[9][11];
assign L2[10][11] = L1[10][11];
assign L2[11][11] = L1[11][11];

assign L2[0][12] = L1[0][12];
assign L2[1][12] = L1[1][12];
assign L2[2][12] = L1[2][12];
assign L2[3][12] = L1[3][12];
assign L2[4][12] = L1[4][12];
assign L2[5][12] = L1[5][12];
assign L2[6][12] = L1[6][12];
assign L2[7][12] = L1[7][12];
assign L2[8][12] = L1[8][12];
assign L2[9][12] = L1[9][12];
assign L2[10][12] = L1[10][12];
assign L2[11][12] = L1[11][12];
assign L2[12][12] = L1[12][12];

assign { L2[0][13+1], L2[0][13] } = L1[0][13] + L1[0+1][13];
assign L2[1][13] = L1[2][13];
assign L2[2][13] = L1[3][13];
assign L2[3][13] = L1[4][13];
assign L2[4][13] = L1[5][13];
assign L2[5][13] = L1[6][13];
assign L2[6][13] = L1[7][13];
assign L2[7][13] = L1[8][13];
assign L2[8][13] = L1[9][13];
assign L2[9][13] = L1[10][13];
assign L2[10][13] = L1[11][13];
assign L2[11][13] = L1[12][13];
assign L2[12][13] = L1[13][13];

assign { L2[0][14+1], L2[1][14] } = L1[0][14] + L1[0+1][14] + L1[0+2][14];
assign { L2[1][14+1], L2[2][14] } = L1[3][14] + L1[3+1][14];
assign L2[3][14] = L1[5][14];
assign L2[4][14] = L1[6][14];
assign L2[5][14] = L1[7][14];
assign L2[6][14] = L1[8][14];
assign L2[7][14] = L1[9][14];
assign L2[8][14] = L1[10][14];
assign L2[9][14] = L1[11][14];
assign L2[10][14] = L1[12][14];
assign L2[11][14] = L1[13][14];
assign L2[12][14] = L1[14][14];

assign { L2[0][15+1], L2[2][15] } = L1[0][15] + L1[0+1][15] + L1[0+2][15];
assign { L2[1][15+1], L2[3][15] } = L1[3][15] + L1[3+1][15] + L1[3+2][15];
assign { L2[2][15+1], L2[4][15] } = L1[6][15] + L1[6+1][15];
assign L2[5][15] = L1[8][15];
assign L2[6][15] = L1[9][15];
assign L2[7][15] = L1[10][15];
assign L2[8][15] = L1[11][15];
assign L2[9][15] = L1[12][15];
assign L2[10][15] = L1[13][15];
assign L2[11][15] = L1[14][15];
assign L2[12][15] = L1[15][15];

assign { L2[0][16+1], L2[3][16] } = L1[0][16] + L1[0+1][16] + L1[0+2][16];
assign { L2[1][16+1], L2[4][16] } = L1[3][16] + L1[3+1][16] + L1[3+2][16];
assign { L2[2][16+1], L2[5][16] } = L1[6][16] + L1[6+1][16] + L1[6+2][16];
assign { L2[3][16+1], L2[6][16] } = L1[9][16] + L1[9+1][16];
assign L2[7][16] = L1[11][16];
assign L2[8][16] = L1[12][16];
assign L2[9][16] = L1[13][16];
assign L2[10][16] = L1[14][16];
assign L2[11][16] = L1[15][16];
assign L2[12][16] = L1[16][16];

assign { L2[0][17+1], L2[4][17] } = L1[0][17] + L1[0+1][17] + L1[0+2][17];
assign { L2[1][17+1], L2[5][17] } = L1[3][17] + L1[3+1][17] + L1[3+2][17];
assign { L2[2][17+1], L2[6][17] } = L1[6][17] + L1[6+1][17] + L1[6+2][17];
assign { L2[3][17+1], L2[7][17] } = L1[9][17] + L1[9+1][17] + L1[9+2][17];
assign { L2[4][17+1], L2[8][17] } = L1[12][17] + L1[12+1][17];
assign L2[9][17] = L1[14][17];
assign L2[10][17] = L1[15][17];
assign L2[11][17] = L1[16][17];
assign L2[12][17] = L1[17][17];

assign { L2[0][18+1], L2[5][18] } = L1[0][18] + L1[0+1][18] + L1[0+2][18];
assign { L2[1][18+1], L2[6][18] } = L1[3][18] + L1[3+1][18] + L1[3+2][18];
assign { L2[2][18+1], L2[7][18] } = L1[6][18] + L1[6+1][18] + L1[6+2][18];
assign { L2[3][18+1], L2[8][18] } = L1[9][18] + L1[9+1][18] + L1[9+2][18];
assign { L2[4][18+1], L2[9][18] } = L1[12][18] + L1[12+1][18] + L1[12+2][18];
assign { L2[5][18+1], L2[10][18] } = L1[15][18] + L1[15+1][18];
assign L2[11][18] = L1[17][18];
assign L2[12][18] = L1[18][18];

assign { L2[0][19+1], L2[6][19] } = L1[0][19] + L1[0+1][19] + L1[0+2][19];
assign { L2[1][19+1], L2[7][19] } = L1[3][19] + L1[3+1][19] + L1[3+2][19];
assign { L2[2][19+1], L2[8][19] } = L1[6][19] + L1[6+1][19] + L1[6+2][19];
assign { L2[3][19+1], L2[9][19] } = L1[9][19] + L1[9+1][19] + L1[9+2][19];
assign { L2[4][19+1], L2[10][19] } = L1[12][19] + L1[12+1][19] + L1[12+2][19];
assign { L2[5][19+1], L2[11][19] } = L1[15][19] + L1[15+1][19] + L1[15+2][19];
assign L2[12][19] = L1[18][19];

assign { L2[0][20+1], L2[6][20] } = L1[0][20] + L1[0+1][20] + L1[0+2][20];
assign { L2[1][20+1], L2[7][20] } = L1[3][20] + L1[3+1][20] + L1[3+2][20];
assign { L2[2][20+1], L2[8][20] } = L1[6][20] + L1[6+1][20] + L1[6+2][20];
assign { L2[3][20+1], L2[9][20] } = L1[9][20] + L1[9+1][20] + L1[9+2][20];
assign { L2[4][20+1], L2[10][20] } = L1[12][20] + L1[12+1][20] + L1[12+2][20];
assign { L2[5][20+1], L2[11][20] } = L1[15][20] + L1[15+1][20] + L1[15+2][20];
assign L2[12][20] = L1[18][20];

assign { L2[0][21+1], L2[6][21] } = L1[0][21] + L1[0+1][21] + L1[0+2][21];
assign { L2[1][21+1], L2[7][21] } = L1[3][21] + L1[3+1][21] + L1[3+2][21];
assign { L2[2][21+1], L2[8][21] } = L1[6][21] + L1[6+1][21] + L1[6+2][21];
assign { L2[3][21+1], L2[9][21] } = L1[9][21] + L1[9+1][21] + L1[9+2][21];
assign { L2[4][21+1], L2[10][21] } = L1[12][21] + L1[12+1][21] + L1[12+2][21];
assign { L2[5][21+1], L2[11][21] } = L1[15][21] + L1[15+1][21] + L1[15+2][21];
assign L2[12][21] = L1[18][21];

assign { L2[0][22+1], L2[6][22] } = L1[0][22] + L1[0+1][22] + L1[0+2][22];
assign { L2[1][22+1], L2[7][22] } = L1[3][22] + L1[3+1][22] + L1[3+2][22];
assign { L2[2][22+1], L2[8][22] } = L1[6][22] + L1[6+1][22] + L1[6+2][22];
assign { L2[3][22+1], L2[9][22] } = L1[9][22] + L1[9+1][22] + L1[9+2][22];
assign { L2[4][22+1], L2[10][22] } = L1[12][22] + L1[12+1][22] + L1[12+2][22];
assign { L2[5][22+1], L2[11][22] } = L1[15][22] + L1[15+1][22] + L1[15+2][22];
assign L2[12][22] = L1[18][22];

assign { L2[0][23+1], L2[6][23] } = L1[0][23] + L1[0+1][23] + L1[0+2][23];
assign { L2[1][23+1], L2[7][23] } = L1[3][23] + L1[3+1][23] + L1[3+2][23];
assign { L2[2][23+1], L2[8][23] } = L1[6][23] + L1[6+1][23] + L1[6+2][23];
assign { L2[3][23+1], L2[9][23] } = L1[9][23] + L1[9+1][23] + L1[9+2][23];
assign { L2[4][23+1], L2[10][23] } = L1[12][23] + L1[12+1][23] + L1[12+2][23];
assign { L2[5][23+1], L2[11][23] } = L1[15][23] + L1[15+1][23] + L1[15+2][23];
assign L2[12][23] = L1[18][23];

assign { L2[0][24+1], L2[6][24] } = L1[0][24] + L1[0+1][24] + L1[0+2][24];
assign { L2[1][24+1], L2[7][24] } = L1[3][24] + L1[3+1][24] + L1[3+2][24];
assign { L2[2][24+1], L2[8][24] } = L1[6][24] + L1[6+1][24] + L1[6+2][24];
assign { L2[3][24+1], L2[9][24] } = L1[9][24] + L1[9+1][24] + L1[9+2][24];
assign { L2[4][24+1], L2[10][24] } = L1[12][24] + L1[12+1][24] + L1[12+2][24];
assign { L2[5][24+1], L2[11][24] } = L1[15][24] + L1[15+1][24] + L1[15+2][24];
assign L2[12][24] = L1[18][24];

assign { L2[0][25+1], L2[6][25] } = L1[0][25] + L1[0+1][25] + L1[0+2][25];
assign { L2[1][25+1], L2[7][25] } = L1[3][25] + L1[3+1][25] + L1[3+2][25];
assign { L2[2][25+1], L2[8][25] } = L1[6][25] + L1[6+1][25] + L1[6+2][25];
assign { L2[3][25+1], L2[9][25] } = L1[9][25] + L1[9+1][25] + L1[9+2][25];
assign { L2[4][25+1], L2[10][25] } = L1[12][25] + L1[12+1][25] + L1[12+2][25];
assign { L2[5][25+1], L2[11][25] } = L1[15][25] + L1[15+1][25] + L1[15+2][25];
assign L2[12][25] = L1[18][25];

assign { L2[0][26+1], L2[6][26] } = L1[0][26] + L1[0+1][26] + L1[0+2][26];
assign { L2[1][26+1], L2[7][26] } = L1[3][26] + L1[3+1][26] + L1[3+2][26];
assign { L2[2][26+1], L2[8][26] } = L1[6][26] + L1[6+1][26] + L1[6+2][26];
assign { L2[3][26+1], L2[9][26] } = L1[9][26] + L1[9+1][26] + L1[9+2][26];
assign { L2[4][26+1], L2[10][26] } = L1[12][26] + L1[12+1][26] + L1[12+2][26];
assign { L2[5][26+1], L2[11][26] } = L1[15][26] + L1[15+1][26] + L1[15+2][26];
assign L2[12][26] = L1[18][26];

assign { L2[0][27+1], L2[6][27] } = L1[0][27] + L1[0+1][27] + L1[0+2][27];
assign { L2[1][27+1], L2[7][27] } = L1[3][27] + L1[3+1][27] + L1[3+2][27];
assign { L2[2][27+1], L2[8][27] } = L1[6][27] + L1[6+1][27] + L1[6+2][27];
assign { L2[3][27+1], L2[9][27] } = L1[9][27] + L1[9+1][27] + L1[9+2][27];
assign { L2[4][27+1], L2[10][27] } = L1[12][27] + L1[12+1][27] + L1[12+2][27];
assign { L2[5][27+1], L2[11][27] } = L1[15][27] + L1[15+1][27] + L1[15+2][27];
assign L2[12][27] = L1[18][27];

assign { L2[0][28+1], L2[6][28] } = L1[0][28] + L1[0+1][28] + L1[0+2][28];
assign { L2[1][28+1], L2[7][28] } = L1[3][28] + L1[3+1][28] + L1[3+2][28];
assign { L2[2][28+1], L2[8][28] } = L1[6][28] + L1[6+1][28] + L1[6+2][28];
assign { L2[3][28+1], L2[9][28] } = L1[9][28] + L1[9+1][28] + L1[9+2][28];
assign { L2[4][28+1], L2[10][28] } = L1[12][28] + L1[12+1][28] + L1[12+2][28];
assign { L2[5][28+1], L2[11][28] } = L1[15][28] + L1[15+1][28] + L1[15+2][28];
assign L2[12][28] = L1[18][28];

assign { L2[0][29+1], L2[6][29] } = L1[0][29] + L1[0+1][29] + L1[0+2][29];
assign { L2[1][29+1], L2[7][29] } = L1[3][29] + L1[3+1][29] + L1[3+2][29];
assign { L2[2][29+1], L2[8][29] } = L1[6][29] + L1[6+1][29] + L1[6+2][29];
assign { L2[3][29+1], L2[9][29] } = L1[9][29] + L1[9+1][29] + L1[9+2][29];
assign { L2[4][29+1], L2[10][29] } = L1[12][29] + L1[12+1][29] + L1[12+2][29];
assign { L2[5][29+1], L2[11][29] } = L1[15][29] + L1[15+1][29] + L1[15+2][29];
assign L2[12][29] = L1[18][29];

assign { L2[0][30+1], L2[6][30] } = L1[0][30] + L1[0+1][30] + L1[0+2][30];
assign { L2[1][30+1], L2[7][30] } = L1[3][30] + L1[3+1][30] + L1[3+2][30];
assign { L2[2][30+1], L2[8][30] } = L1[6][30] + L1[6+1][30] + L1[6+2][30];
assign { L2[3][30+1], L2[9][30] } = L1[9][30] + L1[9+1][30] + L1[9+2][30];
assign { L2[4][30+1], L2[10][30] } = L1[12][30] + L1[12+1][30] + L1[12+2][30];
assign L2[11][30] = L1[15][30];
assign L2[12][30] = L1[16][30];

assign { L2[0][31+1], L2[5][31] } = L1[0][31] + L1[0+1][31] + L1[0+2][31];
assign { L2[1][31+1], L2[6][31] } = L1[3][31] + L1[3+1][31] + L1[3+2][31];
assign { L2[2][31+1], L2[7][31] } = L1[6][31] + L1[6+1][31] + L1[6+2][31];
assign { L2[3][31+1], L2[8][31] } = L1[9][31] + L1[9+1][31] + L1[9+2][31];
assign L2[9][31] = L1[12][31];
assign L2[10][31] = L1[13][31];
assign L2[11][31] = L1[14][31];
assign L2[12][31] = L1[15][31];

assign { L2[0][32+1], L2[4][32] } = L1[0][32] + L1[0+1][32] + L1[0+2][32];
assign { L2[1][32+1], L2[5][32] } = L1[3][32] + L1[3+1][32] + L1[3+2][32];
assign { L2[2][32+1], L2[6][32] } = L1[6][32] + L1[6+1][32] + L1[6+2][32];
assign L2[7][32] = L1[9][32];
assign L2[8][32] = L1[10][32];
assign L2[9][32] = L1[11][32];
assign L2[10][32] = L1[12][32];
assign L2[11][32] = L1[13][32];
assign L2[12][32] = L1[14][32];

assign { L2[0][33+1], L2[3][33] } = L1[0][33] + L1[0+1][33] + L1[0+2][33];
assign { L2[1][33+1], L2[4][33] } = L1[3][33] + L1[3+1][33] + L1[3+2][33];
assign L2[5][33] = L1[6][33];
assign L2[6][33] = L1[7][33];
assign L2[7][33] = L1[8][33];
assign L2[8][33] = L1[9][33];
assign L2[9][33] = L1[10][33];
assign L2[10][33] = L1[11][33];
assign L2[11][33] = L1[12][33];
assign L2[12][33] = L1[13][33];

assign { L2[0][34+1], L2[2][34] } = L1[0][34] + L1[0+1][34] + L1[0+2][34];
assign L2[3][34] = L1[3][34];
assign L2[4][34] = L1[4][34];
assign L2[5][34] = L1[5][34];
assign L2[6][34] = L1[6][34];
assign L2[7][34] = L1[7][34];
assign L2[8][34] = L1[8][34];
assign L2[9][34] = L1[9][34];
assign L2[10][34] = L1[10][34];
assign L2[11][34] = L1[11][34];
assign L2[12][34] = L1[12][34];

assign L2[1][35] = L1[0][35];
assign L2[2][35] = L1[1][35];
assign L2[3][35] = L1[2][35];
assign L2[4][35] = L1[3][35];
assign L2[5][35] = L1[4][35];
assign L2[6][35] = L1[5][35];
assign L2[7][35] = L1[6][35];
assign L2[8][35] = L1[7][35];
assign L2[9][35] = L1[8][35];
assign L2[10][35] = L1[9][35];
assign L2[11][35] = L1[10][35];
assign L2[12][35] = L1[11][35];

assign L2[0][36] = L1[0][36];
assign L2[1][36] = L1[1][36];
assign L2[2][36] = L1[2][36];
assign L2[3][36] = L1[3][36];
assign L2[4][36] = L1[4][36];
assign L2[5][36] = L1[5][36];
assign L2[6][36] = L1[6][36];
assign L2[7][36] = L1[7][36];
assign L2[8][36] = L1[8][36];
assign L2[9][36] = L1[9][36];
assign L2[10][36] = L1[10][36];

assign L2[0][37] = L1[0][37];
assign L2[1][37] = L1[1][37];
assign L2[2][37] = L1[2][37];
assign L2[3][37] = L1[3][37];
assign L2[4][37] = L1[4][37];
assign L2[5][37] = L1[5][37];
assign L2[6][37] = L1[6][37];
assign L2[7][37] = L1[7][37];
assign L2[8][37] = L1[8][37];
assign L2[9][37] = L1[9][37];

assign L2[0][38] = L1[0][38];
assign L2[1][38] = L1[1][38];
assign L2[2][38] = L1[2][38];
assign L2[3][38] = L1[3][38];
assign L2[4][38] = L1[4][38];
assign L2[5][38] = L1[5][38];
assign L2[6][38] = L1[6][38];
assign L2[7][38] = L1[7][38];
assign L2[8][38] = L1[8][38];

assign L2[0][39] = L1[0][39];
assign L2[1][39] = L1[1][39];
assign L2[2][39] = L1[2][39];
assign L2[3][39] = L1[3][39];
assign L2[4][39] = L1[4][39];
assign L2[5][39] = L1[5][39];
assign L2[6][39] = L1[6][39];
assign L2[7][39] = L1[7][39];

assign L2[0][40] = L1[0][40];
assign L2[1][40] = L1[1][40];
assign L2[2][40] = L1[2][40];
assign L2[3][40] = L1[3][40];
assign L2[4][40] = L1[4][40];
assign L2[5][40] = L1[5][40];
assign L2[6][40] = L1[6][40];

assign L2[0][41] = L1[0][41];
assign L2[1][41] = L1[1][41];
assign L2[2][41] = L1[2][41];
assign L2[3][41] = L1[3][41];
assign L2[4][41] = L1[4][41];
assign L2[5][41] = L1[5][41];

assign L2[0][42] = L1[0][42];
assign L2[1][42] = L1[1][42];
assign L2[2][42] = L1[2][42];
assign L2[3][42] = L1[3][42];
assign L2[4][42] = L1[4][42];

assign L2[0][43] = L1[0][43];
assign L2[1][43] = L1[1][43];
assign L2[2][43] = L1[2][43];
assign L2[3][43] = L1[3][43];

assign L2[0][44] = L1[0][44];
assign L2[1][44] = L1[1][44];
assign L2[2][44] = L1[2][44];

assign L2[0][45] = L1[0][45];
assign L2[1][45] = L1[1][45];

assign L2[0][46] = L1[0][46];


assign L3[0][0] = L2[0][0];

assign L3[0][1] = L2[0][1];
assign L3[1][1] = L2[1][1];

assign L3[0][2] = L2[0][2];
assign L3[1][2] = L2[1][2];
assign L3[2][2] = L2[2][2];

assign L3[0][3] = L2[0][3];
assign L3[1][3] = L2[1][3];
assign L3[2][3] = L2[2][3];
assign L3[3][3] = L2[3][3];

assign L3[0][4] = L2[0][4];
assign L3[1][4] = L2[1][4];
assign L3[2][4] = L2[2][4];
assign L3[3][4] = L2[3][4];
assign L3[4][4] = L2[4][4];

assign L3[0][5] = L2[0][5];
assign L3[1][5] = L2[1][5];
assign L3[2][5] = L2[2][5];
assign L3[3][5] = L2[3][5];
assign L3[4][5] = L2[4][5];
assign L3[5][5] = L2[5][5];

assign L3[0][6] = L2[0][6];
assign L3[1][6] = L2[1][6];
assign L3[2][6] = L2[2][6];
assign L3[3][6] = L2[3][6];
assign L3[4][6] = L2[4][6];
assign L3[5][6] = L2[5][6];
assign L3[6][6] = L2[6][6];

assign L3[0][7] = L2[0][7];
assign L3[1][7] = L2[1][7];
assign L3[2][7] = L2[2][7];
assign L3[3][7] = L2[3][7];
assign L3[4][7] = L2[4][7];
assign L3[5][7] = L2[5][7];
assign L3[6][7] = L2[6][7];
assign L3[7][7] = L2[7][7];

assign L3[0][8] = L2[0][8];
assign L3[1][8] = L2[1][8];
assign L3[2][8] = L2[2][8];
assign L3[3][8] = L2[3][8];
assign L3[4][8] = L2[4][8];
assign L3[5][8] = L2[5][8];
assign L3[6][8] = L2[6][8];
assign L3[7][8] = L2[7][8];
assign L3[8][8] = L2[8][8];

assign { L3[0][9+1], L3[0][9] } = L2[0][9] + L2[0+1][9];
assign L3[1][9] = L2[2][9];
assign L3[2][9] = L2[3][9];
assign L3[3][9] = L2[4][9];
assign L3[4][9] = L2[5][9];
assign L3[5][9] = L2[6][9];
assign L3[6][9] = L2[7][9];
assign L3[7][9] = L2[8][9];
assign L3[8][9] = L2[9][9];

assign { L3[0][10+1], L3[1][10] } = L2[0][10] + L2[0+1][10] + L2[0+2][10];
assign { L3[1][10+1], L3[2][10] } = L2[3][10] + L2[3+1][10];
assign L3[3][10] = L2[5][10];
assign L3[4][10] = L2[6][10];
assign L3[5][10] = L2[7][10];
assign L3[6][10] = L2[8][10];
assign L3[7][10] = L2[9][10];
assign L3[8][10] = L2[10][10];

assign { L3[0][11+1], L3[2][11] } = L2[0][11] + L2[0+1][11] + L2[0+2][11];
assign { L3[1][11+1], L3[3][11] } = L2[3][11] + L2[3+1][11] + L2[3+2][11];
assign { L3[2][11+1], L3[4][11] } = L2[6][11] + L2[6+1][11];
assign L3[5][11] = L2[8][11];
assign L3[6][11] = L2[9][11];
assign L3[7][11] = L2[10][11];
assign L3[8][11] = L2[11][11];

assign { L3[0][12+1], L3[3][12] } = L2[0][12] + L2[0+1][12] + L2[0+2][12];
assign { L3[1][12+1], L3[4][12] } = L2[3][12] + L2[3+1][12] + L2[3+2][12];
assign { L3[2][12+1], L3[5][12] } = L2[6][12] + L2[6+1][12] + L2[6+2][12];
assign { L3[3][12+1], L3[6][12] } = L2[9][12] + L2[9+1][12];
assign L3[7][12] = L2[11][12];
assign L3[8][12] = L2[12][12];

assign { L3[0][13+1], L3[4][13] } = L2[0][13] + L2[0+1][13] + L2[0+2][13];
assign { L3[1][13+1], L3[5][13] } = L2[3][13] + L2[3+1][13] + L2[3+2][13];
assign { L3[2][13+1], L3[6][13] } = L2[6][13] + L2[6+1][13] + L2[6+2][13];
assign { L3[3][13+1], L3[7][13] } = L2[9][13] + L2[9+1][13] + L2[9+2][13];
assign L3[8][13] = L2[12][13];

assign { L3[0][14+1], L3[4][14] } = L2[0][14] + L2[0+1][14] + L2[0+2][14];
assign { L3[1][14+1], L3[5][14] } = L2[3][14] + L2[3+1][14] + L2[3+2][14];
assign { L3[2][14+1], L3[6][14] } = L2[6][14] + L2[6+1][14] + L2[6+2][14];
assign { L3[3][14+1], L3[7][14] } = L2[9][14] + L2[9+1][14] + L2[9+2][14];
assign L3[8][14] = L2[12][14];

assign { L3[0][15+1], L3[4][15] } = L2[0][15] + L2[0+1][15] + L2[0+2][15];
assign { L3[1][15+1], L3[5][15] } = L2[3][15] + L2[3+1][15] + L2[3+2][15];
assign { L3[2][15+1], L3[6][15] } = L2[6][15] + L2[6+1][15] + L2[6+2][15];
assign { L3[3][15+1], L3[7][15] } = L2[9][15] + L2[9+1][15] + L2[9+2][15];
assign L3[8][15] = L2[12][15];

assign { L3[0][16+1], L3[4][16] } = L2[0][16] + L2[0+1][16] + L2[0+2][16];
assign { L3[1][16+1], L3[5][16] } = L2[3][16] + L2[3+1][16] + L2[3+2][16];
assign { L3[2][16+1], L3[6][16] } = L2[6][16] + L2[6+1][16] + L2[6+2][16];
assign { L3[3][16+1], L3[7][16] } = L2[9][16] + L2[9+1][16] + L2[9+2][16];
assign L3[8][16] = L2[12][16];

assign { L3[0][17+1], L3[4][17] } = L2[0][17] + L2[0+1][17] + L2[0+2][17];
assign { L3[1][17+1], L3[5][17] } = L2[3][17] + L2[3+1][17] + L2[3+2][17];
assign { L3[2][17+1], L3[6][17] } = L2[6][17] + L2[6+1][17] + L2[6+2][17];
assign { L3[3][17+1], L3[7][17] } = L2[9][17] + L2[9+1][17] + L2[9+2][17];
assign L3[8][17] = L2[12][17];

assign { L3[0][18+1], L3[4][18] } = L2[0][18] + L2[0+1][18] + L2[0+2][18];
assign { L3[1][18+1], L3[5][18] } = L2[3][18] + L2[3+1][18] + L2[3+2][18];
assign { L3[2][18+1], L3[6][18] } = L2[6][18] + L2[6+1][18] + L2[6+2][18];
assign { L3[3][18+1], L3[7][18] } = L2[9][18] + L2[9+1][18] + L2[9+2][18];
assign L3[8][18] = L2[12][18];

assign { L3[0][19+1], L3[4][19] } = L2[0][19] + L2[0+1][19] + L2[0+2][19];
assign { L3[1][19+1], L3[5][19] } = L2[3][19] + L2[3+1][19] + L2[3+2][19];
assign { L3[2][19+1], L3[6][19] } = L2[6][19] + L2[6+1][19] + L2[6+2][19];
assign { L3[3][19+1], L3[7][19] } = L2[9][19] + L2[9+1][19] + L2[9+2][19];
assign L3[8][19] = L2[12][19];

assign { L3[0][20+1], L3[4][20] } = L2[0][20] + L2[0+1][20] + L2[0+2][20];
assign { L3[1][20+1], L3[5][20] } = L2[3][20] + L2[3+1][20] + L2[3+2][20];
assign { L3[2][20+1], L3[6][20] } = L2[6][20] + L2[6+1][20] + L2[6+2][20];
assign { L3[3][20+1], L3[7][20] } = L2[9][20] + L2[9+1][20] + L2[9+2][20];
assign L3[8][20] = L2[12][20];

assign { L3[0][21+1], L3[4][21] } = L2[0][21] + L2[0+1][21] + L2[0+2][21];
assign { L3[1][21+1], L3[5][21] } = L2[3][21] + L2[3+1][21] + L2[3+2][21];
assign { L3[2][21+1], L3[6][21] } = L2[6][21] + L2[6+1][21] + L2[6+2][21];
assign { L3[3][21+1], L3[7][21] } = L2[9][21] + L2[9+1][21] + L2[9+2][21];
assign L3[8][21] = L2[12][21];

assign { L3[0][22+1], L3[4][22] } = L2[0][22] + L2[0+1][22] + L2[0+2][22];
assign { L3[1][22+1], L3[5][22] } = L2[3][22] + L2[3+1][22] + L2[3+2][22];
assign { L3[2][22+1], L3[6][22] } = L2[6][22] + L2[6+1][22] + L2[6+2][22];
assign { L3[3][22+1], L3[7][22] } = L2[9][22] + L2[9+1][22] + L2[9+2][22];
assign L3[8][22] = L2[12][22];

assign { L3[0][23+1], L3[4][23] } = L2[0][23] + L2[0+1][23] + L2[0+2][23];
assign { L3[1][23+1], L3[5][23] } = L2[3][23] + L2[3+1][23] + L2[3+2][23];
assign { L3[2][23+1], L3[6][23] } = L2[6][23] + L2[6+1][23] + L2[6+2][23];
assign { L3[3][23+1], L3[7][23] } = L2[9][23] + L2[9+1][23] + L2[9+2][23];
assign L3[8][23] = L2[12][23];

assign { L3[0][24+1], L3[4][24] } = L2[0][24] + L2[0+1][24] + L2[0+2][24];
assign { L3[1][24+1], L3[5][24] } = L2[3][24] + L2[3+1][24] + L2[3+2][24];
assign { L3[2][24+1], L3[6][24] } = L2[6][24] + L2[6+1][24] + L2[6+2][24];
assign { L3[3][24+1], L3[7][24] } = L2[9][24] + L2[9+1][24] + L2[9+2][24];
assign L3[8][24] = L2[12][24];

assign { L3[0][25+1], L3[4][25] } = L2[0][25] + L2[0+1][25] + L2[0+2][25];
assign { L3[1][25+1], L3[5][25] } = L2[3][25] + L2[3+1][25] + L2[3+2][25];
assign { L3[2][25+1], L3[6][25] } = L2[6][25] + L2[6+1][25] + L2[6+2][25];
assign { L3[3][25+1], L3[7][25] } = L2[9][25] + L2[9+1][25] + L2[9+2][25];
assign L3[8][25] = L2[12][25];

assign { L3[0][26+1], L3[4][26] } = L2[0][26] + L2[0+1][26] + L2[0+2][26];
assign { L3[1][26+1], L3[5][26] } = L2[3][26] + L2[3+1][26] + L2[3+2][26];
assign { L3[2][26+1], L3[6][26] } = L2[6][26] + L2[6+1][26] + L2[6+2][26];
assign { L3[3][26+1], L3[7][26] } = L2[9][26] + L2[9+1][26] + L2[9+2][26];
assign L3[8][26] = L2[12][26];

assign { L3[0][27+1], L3[4][27] } = L2[0][27] + L2[0+1][27] + L2[0+2][27];
assign { L3[1][27+1], L3[5][27] } = L2[3][27] + L2[3+1][27] + L2[3+2][27];
assign { L3[2][27+1], L3[6][27] } = L2[6][27] + L2[6+1][27] + L2[6+2][27];
assign { L3[3][27+1], L3[7][27] } = L2[9][27] + L2[9+1][27] + L2[9+2][27];
assign L3[8][27] = L2[12][27];

assign { L3[0][28+1], L3[4][28] } = L2[0][28] + L2[0+1][28] + L2[0+2][28];
assign { L3[1][28+1], L3[5][28] } = L2[3][28] + L2[3+1][28] + L2[3+2][28];
assign { L3[2][28+1], L3[6][28] } = L2[6][28] + L2[6+1][28] + L2[6+2][28];
assign { L3[3][28+1], L3[7][28] } = L2[9][28] + L2[9+1][28] + L2[9+2][28];
assign L3[8][28] = L2[12][28];

assign { L3[0][29+1], L3[4][29] } = L2[0][29] + L2[0+1][29] + L2[0+2][29];
assign { L3[1][29+1], L3[5][29] } = L2[3][29] + L2[3+1][29] + L2[3+2][29];
assign { L3[2][29+1], L3[6][29] } = L2[6][29] + L2[6+1][29] + L2[6+2][29];
assign { L3[3][29+1], L3[7][29] } = L2[9][29] + L2[9+1][29] + L2[9+2][29];
assign L3[8][29] = L2[12][29];

assign { L3[0][30+1], L3[4][30] } = L2[0][30] + L2[0+1][30] + L2[0+2][30];
assign { L3[1][30+1], L3[5][30] } = L2[3][30] + L2[3+1][30] + L2[3+2][30];
assign { L3[2][30+1], L3[6][30] } = L2[6][30] + L2[6+1][30] + L2[6+2][30];
assign { L3[3][30+1], L3[7][30] } = L2[9][30] + L2[9+1][30] + L2[9+2][30];
assign L3[8][30] = L2[12][30];

assign { L3[0][31+1], L3[4][31] } = L2[0][31] + L2[0+1][31] + L2[0+2][31];
assign { L3[1][31+1], L3[5][31] } = L2[3][31] + L2[3+1][31] + L2[3+2][31];
assign { L3[2][31+1], L3[6][31] } = L2[6][31] + L2[6+1][31] + L2[6+2][31];
assign { L3[3][31+1], L3[7][31] } = L2[9][31] + L2[9+1][31] + L2[9+2][31];
assign L3[8][31] = L2[12][31];

assign { L3[0][32+1], L3[4][32] } = L2[0][32] + L2[0+1][32] + L2[0+2][32];
assign { L3[1][32+1], L3[5][32] } = L2[3][32] + L2[3+1][32] + L2[3+2][32];
assign { L3[2][32+1], L3[6][32] } = L2[6][32] + L2[6+1][32] + L2[6+2][32];
assign { L3[3][32+1], L3[7][32] } = L2[9][32] + L2[9+1][32] + L2[9+2][32];
assign L3[8][32] = L2[12][32];

assign { L3[0][33+1], L3[4][33] } = L2[0][33] + L2[0+1][33] + L2[0+2][33];
assign { L3[1][33+1], L3[5][33] } = L2[3][33] + L2[3+1][33] + L2[3+2][33];
assign { L3[2][33+1], L3[6][33] } = L2[6][33] + L2[6+1][33] + L2[6+2][33];
assign { L3[3][33+1], L3[7][33] } = L2[9][33] + L2[9+1][33] + L2[9+2][33];
assign L3[8][33] = L2[12][33];

assign { L3[0][34+1], L3[4][34] } = L2[0][34] + L2[0+1][34] + L2[0+2][34];
assign { L3[1][34+1], L3[5][34] } = L2[3][34] + L2[3+1][34] + L2[3+2][34];
assign { L3[2][34+1], L3[6][34] } = L2[6][34] + L2[6+1][34] + L2[6+2][34];
assign { L3[3][34+1], L3[7][34] } = L2[9][34] + L2[9+1][34] + L2[9+2][34];
assign L3[8][34] = L2[12][34];

assign { L3[0][35+1], L3[4][35] } = L2[0][35] + L2[0+1][35] + L2[0+2][35];
assign { L3[1][35+1], L3[5][35] } = L2[3][35] + L2[3+1][35] + L2[3+2][35];
assign { L3[2][35+1], L3[6][35] } = L2[6][35] + L2[6+1][35] + L2[6+2][35];
assign { L3[3][35+1], L3[7][35] } = L2[9][35] + L2[9+1][35] + L2[9+2][35];
assign L3[8][35] = L2[12][35];

assign { L3[0][36+1], L3[4][36] } = L2[0][36] + L2[0+1][36] + L2[0+2][36];
assign { L3[1][36+1], L3[5][36] } = L2[3][36] + L2[3+1][36] + L2[3+2][36];
assign { L3[2][36+1], L3[6][36] } = L2[6][36] + L2[6+1][36] + L2[6+2][36];
assign L3[7][36] = L2[9][36];
assign L3[8][36] = L2[10][36];

assign { L3[0][37+1], L3[3][37] } = L2[0][37] + L2[0+1][37] + L2[0+2][37];
assign { L3[1][37+1], L3[4][37] } = L2[3][37] + L2[3+1][37] + L2[3+2][37];
assign L3[5][37] = L2[6][37];
assign L3[6][37] = L2[7][37];
assign L3[7][37] = L2[8][37];
assign L3[8][37] = L2[9][37];

assign { L3[0][38+1], L3[2][38] } = L2[0][38] + L2[0+1][38] + L2[0+2][38];
assign L3[3][38] = L2[3][38];
assign L3[4][38] = L2[4][38];
assign L3[5][38] = L2[5][38];
assign L3[6][38] = L2[6][38];
assign L3[7][38] = L2[7][38];
assign L3[8][38] = L2[8][38];

assign L3[1][39] = L2[0][39];
assign L3[2][39] = L2[1][39];
assign L3[3][39] = L2[2][39];
assign L3[4][39] = L2[3][39];
assign L3[5][39] = L2[4][39];
assign L3[6][39] = L2[5][39];
assign L3[7][39] = L2[6][39];
assign L3[8][39] = L2[7][39];

assign L3[0][40] = L2[0][40];
assign L3[1][40] = L2[1][40];
assign L3[2][40] = L2[2][40];
assign L3[3][40] = L2[3][40];
assign L3[4][40] = L2[4][40];
assign L3[5][40] = L2[5][40];
assign L3[6][40] = L2[6][40];

assign L3[0][41] = L2[0][41];
assign L3[1][41] = L2[1][41];
assign L3[2][41] = L2[2][41];
assign L3[3][41] = L2[3][41];
assign L3[4][41] = L2[4][41];
assign L3[5][41] = L2[5][41];

assign L3[0][42] = L2[0][42];
assign L3[1][42] = L2[1][42];
assign L3[2][42] = L2[2][42];
assign L3[3][42] = L2[3][42];
assign L3[4][42] = L2[4][42];

assign L3[0][43] = L2[0][43];
assign L3[1][43] = L2[1][43];
assign L3[2][43] = L2[2][43];
assign L3[3][43] = L2[3][43];

assign L3[0][44] = L2[0][44];
assign L3[1][44] = L2[1][44];
assign L3[2][44] = L2[2][44];

assign L3[0][45] = L2[0][45];
assign L3[1][45] = L2[1][45];

assign L3[0][46] = L2[0][46];


assign L4[0][0] = L3[0][0];

assign L4[0][1] = L3[0][1];
assign L4[1][1] = L3[1][1];

assign L4[0][2] = L3[0][2];
assign L4[1][2] = L3[1][2];
assign L4[2][2] = L3[2][2];

assign L4[0][3] = L3[0][3];
assign L4[1][3] = L3[1][3];
assign L4[2][3] = L3[2][3];
assign L4[3][3] = L3[3][3];

assign L4[0][4] = L3[0][4];
assign L4[1][4] = L3[1][4];
assign L4[2][4] = L3[2][4];
assign L4[3][4] = L3[3][4];
assign L4[4][4] = L3[4][4];

assign L4[0][5] = L3[0][5];
assign L4[1][5] = L3[1][5];
assign L4[2][5] = L3[2][5];
assign L4[3][5] = L3[3][5];
assign L4[4][5] = L3[4][5];
assign L4[5][5] = L3[5][5];

assign { L4[0][6+1], L4[0][6] } = L3[0][6] + L3[0+1][6];
assign L4[1][6] = L3[2][6];
assign L4[2][6] = L3[3][6];
assign L4[3][6] = L3[4][6];
assign L4[4][6] = L3[5][6];
assign L4[5][6] = L3[6][6];

assign { L4[0][7+1], L4[1][7] } = L3[0][7] + L3[0+1][7] + L3[0+2][7];
assign { L4[1][7+1], L4[2][7] } = L3[3][7] + L3[3+1][7];
assign L4[3][7] = L3[5][7];
assign L4[4][7] = L3[6][7];
assign L4[5][7] = L3[7][7];

assign { L4[0][8+1], L4[2][8] } = L3[0][8] + L3[0+1][8] + L3[0+2][8];
assign { L4[1][8+1], L4[3][8] } = L3[3][8] + L3[3+1][8] + L3[3+2][8];
assign { L4[2][8+1], L4[4][8] } = L3[6][8] + L3[6+1][8];
assign L4[5][8] = L3[8][8];

assign { L4[0][9+1], L4[3][9] } = L3[0][9] + L3[0+1][9] + L3[0+2][9];
assign { L4[1][9+1], L4[4][9] } = L3[3][9] + L3[3+1][9] + L3[3+2][9];
assign { L4[2][9+1], L4[5][9] } = L3[6][9] + L3[6+1][9] + L3[6+2][9];

assign { L4[0][10+1], L4[3][10] } = L3[0][10] + L3[0+1][10] + L3[0+2][10];
assign { L4[1][10+1], L4[4][10] } = L3[3][10] + L3[3+1][10] + L3[3+2][10];
assign { L4[2][10+1], L4[5][10] } = L3[6][10] + L3[6+1][10] + L3[6+2][10];

assign { L4[0][11+1], L4[3][11] } = L3[0][11] + L3[0+1][11] + L3[0+2][11];
assign { L4[1][11+1], L4[4][11] } = L3[3][11] + L3[3+1][11] + L3[3+2][11];
assign { L4[2][11+1], L4[5][11] } = L3[6][11] + L3[6+1][11] + L3[6+2][11];

assign { L4[0][12+1], L4[3][12] } = L3[0][12] + L3[0+1][12] + L3[0+2][12];
assign { L4[1][12+1], L4[4][12] } = L3[3][12] + L3[3+1][12] + L3[3+2][12];
assign { L4[2][12+1], L4[5][12] } = L3[6][12] + L3[6+1][12] + L3[6+2][12];

assign { L4[0][13+1], L4[3][13] } = L3[0][13] + L3[0+1][13] + L3[0+2][13];
assign { L4[1][13+1], L4[4][13] } = L3[3][13] + L3[3+1][13] + L3[3+2][13];
assign { L4[2][13+1], L4[5][13] } = L3[6][13] + L3[6+1][13] + L3[6+2][13];

assign { L4[0][14+1], L4[3][14] } = L3[0][14] + L3[0+1][14] + L3[0+2][14];
assign { L4[1][14+1], L4[4][14] } = L3[3][14] + L3[3+1][14] + L3[3+2][14];
assign { L4[2][14+1], L4[5][14] } = L3[6][14] + L3[6+1][14] + L3[6+2][14];

assign { L4[0][15+1], L4[3][15] } = L3[0][15] + L3[0+1][15] + L3[0+2][15];
assign { L4[1][15+1], L4[4][15] } = L3[3][15] + L3[3+1][15] + L3[3+2][15];
assign { L4[2][15+1], L4[5][15] } = L3[6][15] + L3[6+1][15] + L3[6+2][15];

assign { L4[0][16+1], L4[3][16] } = L3[0][16] + L3[0+1][16] + L3[0+2][16];
assign { L4[1][16+1], L4[4][16] } = L3[3][16] + L3[3+1][16] + L3[3+2][16];
assign { L4[2][16+1], L4[5][16] } = L3[6][16] + L3[6+1][16] + L3[6+2][16];

assign { L4[0][17+1], L4[3][17] } = L3[0][17] + L3[0+1][17] + L3[0+2][17];
assign { L4[1][17+1], L4[4][17] } = L3[3][17] + L3[3+1][17] + L3[3+2][17];
assign { L4[2][17+1], L4[5][17] } = L3[6][17] + L3[6+1][17] + L3[6+2][17];

assign { L4[0][18+1], L4[3][18] } = L3[0][18] + L3[0+1][18] + L3[0+2][18];
assign { L4[1][18+1], L4[4][18] } = L3[3][18] + L3[3+1][18] + L3[3+2][18];
assign { L4[2][18+1], L4[5][18] } = L3[6][18] + L3[6+1][18] + L3[6+2][18];

assign { L4[0][19+1], L4[3][19] } = L3[0][19] + L3[0+1][19] + L3[0+2][19];
assign { L4[1][19+1], L4[4][19] } = L3[3][19] + L3[3+1][19] + L3[3+2][19];
assign { L4[2][19+1], L4[5][19] } = L3[6][19] + L3[6+1][19] + L3[6+2][19];

assign { L4[0][20+1], L4[3][20] } = L3[0][20] + L3[0+1][20] + L3[0+2][20];
assign { L4[1][20+1], L4[4][20] } = L3[3][20] + L3[3+1][20] + L3[3+2][20];
assign { L4[2][20+1], L4[5][20] } = L3[6][20] + L3[6+1][20] + L3[6+2][20];

assign { L4[0][21+1], L4[3][21] } = L3[0][21] + L3[0+1][21] + L3[0+2][21];
assign { L4[1][21+1], L4[4][21] } = L3[3][21] + L3[3+1][21] + L3[3+2][21];
assign { L4[2][21+1], L4[5][21] } = L3[6][21] + L3[6+1][21] + L3[6+2][21];

assign { L4[0][22+1], L4[3][22] } = L3[0][22] + L3[0+1][22] + L3[0+2][22];
assign { L4[1][22+1], L4[4][22] } = L3[3][22] + L3[3+1][22] + L3[3+2][22];
assign { L4[2][22+1], L4[5][22] } = L3[6][22] + L3[6+1][22] + L3[6+2][22];

assign { L4[0][23+1], L4[3][23] } = L3[0][23] + L3[0+1][23] + L3[0+2][23];
assign { L4[1][23+1], L4[4][23] } = L3[3][23] + L3[3+1][23] + L3[3+2][23];
assign { L4[2][23+1], L4[5][23] } = L3[6][23] + L3[6+1][23] + L3[6+2][23];

assign { L4[0][24+1], L4[3][24] } = L3[0][24] + L3[0+1][24] + L3[0+2][24];
assign { L4[1][24+1], L4[4][24] } = L3[3][24] + L3[3+1][24] + L3[3+2][24];
assign { L4[2][24+1], L4[5][24] } = L3[6][24] + L3[6+1][24] + L3[6+2][24];

assign { L4[0][25+1], L4[3][25] } = L3[0][25] + L3[0+1][25] + L3[0+2][25];
assign { L4[1][25+1], L4[4][25] } = L3[3][25] + L3[3+1][25] + L3[3+2][25];
assign { L4[2][25+1], L4[5][25] } = L3[6][25] + L3[6+1][25] + L3[6+2][25];

assign { L4[0][26+1], L4[3][26] } = L3[0][26] + L3[0+1][26] + L3[0+2][26];
assign { L4[1][26+1], L4[4][26] } = L3[3][26] + L3[3+1][26] + L3[3+2][26];
assign { L4[2][26+1], L4[5][26] } = L3[6][26] + L3[6+1][26] + L3[6+2][26];

assign { L4[0][27+1], L4[3][27] } = L3[0][27] + L3[0+1][27] + L3[0+2][27];
assign { L4[1][27+1], L4[4][27] } = L3[3][27] + L3[3+1][27] + L3[3+2][27];
assign { L4[2][27+1], L4[5][27] } = L3[6][27] + L3[6+1][27] + L3[6+2][27];

assign { L4[0][28+1], L4[3][28] } = L3[0][28] + L3[0+1][28] + L3[0+2][28];
assign { L4[1][28+1], L4[4][28] } = L3[3][28] + L3[3+1][28] + L3[3+2][28];
assign { L4[2][28+1], L4[5][28] } = L3[6][28] + L3[6+1][28] + L3[6+2][28];

assign { L4[0][29+1], L4[3][29] } = L3[0][29] + L3[0+1][29] + L3[0+2][29];
assign { L4[1][29+1], L4[4][29] } = L3[3][29] + L3[3+1][29] + L3[3+2][29];
assign { L4[2][29+1], L4[5][29] } = L3[6][29] + L3[6+1][29] + L3[6+2][29];

assign { L4[0][30+1], L4[3][30] } = L3[0][30] + L3[0+1][30] + L3[0+2][30];
assign { L4[1][30+1], L4[4][30] } = L3[3][30] + L3[3+1][30] + L3[3+2][30];
assign { L4[2][30+1], L4[5][30] } = L3[6][30] + L3[6+1][30] + L3[6+2][30];

assign { L4[0][31+1], L4[3][31] } = L3[0][31] + L3[0+1][31] + L3[0+2][31];
assign { L4[1][31+1], L4[4][31] } = L3[3][31] + L3[3+1][31] + L3[3+2][31];
assign { L4[2][31+1], L4[5][31] } = L3[6][31] + L3[6+1][31] + L3[6+2][31];

assign { L4[0][32+1], L4[3][32] } = L3[0][32] + L3[0+1][32] + L3[0+2][32];
assign { L4[1][32+1], L4[4][32] } = L3[3][32] + L3[3+1][32] + L3[3+2][32];
assign { L4[2][32+1], L4[5][32] } = L3[6][32] + L3[6+1][32] + L3[6+2][32];

assign { L4[0][33+1], L4[3][33] } = L3[0][33] + L3[0+1][33] + L3[0+2][33];
assign { L4[1][33+1], L4[4][33] } = L3[3][33] + L3[3+1][33] + L3[3+2][33];
assign { L4[2][33+1], L4[5][33] } = L3[6][33] + L3[6+1][33] + L3[6+2][33];

assign { L4[0][34+1], L4[3][34] } = L3[0][34] + L3[0+1][34] + L3[0+2][34];
assign { L4[1][34+1], L4[4][34] } = L3[3][34] + L3[3+1][34] + L3[3+2][34];
assign { L4[2][34+1], L4[5][34] } = L3[6][34] + L3[6+1][34] + L3[6+2][34];

assign { L4[0][35+1], L4[3][35] } = L3[0][35] + L3[0+1][35] + L3[0+2][35];
assign { L4[1][35+1], L4[4][35] } = L3[3][35] + L3[3+1][35] + L3[3+2][35];
assign { L4[2][35+1], L4[5][35] } = L3[6][35] + L3[6+1][35] + L3[6+2][35];

assign { L4[0][36+1], L4[3][36] } = L3[0][36] + L3[0+1][36] + L3[0+2][36];
assign { L4[1][36+1], L4[4][36] } = L3[3][36] + L3[3+1][36] + L3[3+2][36];
assign { L4[2][36+1], L4[5][36] } = L3[6][36] + L3[6+1][36] + L3[6+2][36];

assign { L4[0][37+1], L4[3][37] } = L3[0][37] + L3[0+1][37] + L3[0+2][37];
assign { L4[1][37+1], L4[4][37] } = L3[3][37] + L3[3+1][37] + L3[3+2][37];
assign { L4[2][37+1], L4[5][37] } = L3[6][37] + L3[6+1][37] + L3[6+2][37];

assign { L4[0][38+1], L4[3][38] } = L3[0][38] + L3[0+1][38] + L3[0+2][38];
assign { L4[1][38+1], L4[4][38] } = L3[3][38] + L3[3+1][38] + L3[3+2][38];
assign { L4[2][38+1], L4[5][38] } = L3[6][38] + L3[6+1][38] + L3[6+2][38];

assign { L4[0][39+1], L4[3][39] } = L3[0][39] + L3[0+1][39] + L3[0+2][39];
assign { L4[1][39+1], L4[4][39] } = L3[3][39] + L3[3+1][39] + L3[3+2][39];
assign { L4[2][39+1], L4[5][39] } = L3[6][39] + L3[6+1][39] + L3[6+2][39];

assign { L4[0][40+1], L4[3][40] } = L3[0][40] + L3[0+1][40] + L3[0+2][40];
assign { L4[1][40+1], L4[4][40] } = L3[3][40] + L3[3+1][40] + L3[3+2][40];
assign L4[5][40] = L3[6][40];

assign { L4[0][41+1], L4[2][41] } = L3[0][41] + L3[0+1][41] + L3[0+2][41];
assign L4[3][41] = L3[3][41];
assign L4[4][41] = L3[4][41];
assign L4[5][41] = L3[5][41];

assign L4[1][42] = L3[0][42];
assign L4[2][42] = L3[1][42];
assign L4[3][42] = L3[2][42];
assign L4[4][42] = L3[3][42];
assign L4[5][42] = L3[4][42];

assign L4[0][43] = L3[0][43];
assign L4[1][43] = L3[1][43];
assign L4[2][43] = L3[2][43];
assign L4[3][43] = L3[3][43];

assign L4[0][44] = L3[0][44];
assign L4[1][44] = L3[1][44];
assign L4[2][44] = L3[2][44];

assign L4[0][45] = L3[0][45];
assign L4[1][45] = L3[1][45];

assign L4[0][46] = L3[0][46];


assign L5[0][0] = L4[0][0];

assign L5[0][1] = L4[0][1];
assign L5[1][1] = L4[1][1];

assign L5[0][2] = L4[0][2];
assign L5[1][2] = L4[1][2];
assign L5[2][2] = L4[2][2];

assign L5[0][3] = L4[0][3];
assign L5[1][3] = L4[1][3];
assign L5[2][3] = L4[2][3];
assign L5[3][3] = L4[3][3];

assign { L5[0][4+1], L5[0][4] } = L4[0][4] + L4[0+1][4];
assign L5[1][4] = L4[2][4];
assign L5[2][4] = L4[3][4];
assign L5[3][4] = L4[4][4];

assign { L5[0][5+1], L5[1][5] } = L4[0][5] + L4[0+1][5] + L4[0+2][5];
assign { L5[1][5+1], L5[2][5] } = L4[3][5] + L4[3+1][5];
assign L5[3][5] = L4[5][5];

assign { L5[0][6+1], L5[2][6] } = L4[0][6] + L4[0+1][6] + L4[0+2][6];
assign { L5[1][6+1], L5[3][6] } = L4[3][6] + L4[3+1][6] + L4[3+2][6];

assign { L5[0][7+1], L5[2][7] } = L4[0][7] + L4[0+1][7] + L4[0+2][7];
assign { L5[1][7+1], L5[3][7] } = L4[3][7] + L4[3+1][7] + L4[3+2][7];

assign { L5[0][8+1], L5[2][8] } = L4[0][8] + L4[0+1][8] + L4[0+2][8];
assign { L5[1][8+1], L5[3][8] } = L4[3][8] + L4[3+1][8] + L4[3+2][8];

assign { L5[0][9+1], L5[2][9] } = L4[0][9] + L4[0+1][9] + L4[0+2][9];
assign { L5[1][9+1], L5[3][9] } = L4[3][9] + L4[3+1][9] + L4[3+2][9];

assign { L5[0][10+1], L5[2][10] } = L4[0][10] + L4[0+1][10] + L4[0+2][10];
assign { L5[1][10+1], L5[3][10] } = L4[3][10] + L4[3+1][10] + L4[3+2][10];

assign { L5[0][11+1], L5[2][11] } = L4[0][11] + L4[0+1][11] + L4[0+2][11];
assign { L5[1][11+1], L5[3][11] } = L4[3][11] + L4[3+1][11] + L4[3+2][11];

assign { L5[0][12+1], L5[2][12] } = L4[0][12] + L4[0+1][12] + L4[0+2][12];
assign { L5[1][12+1], L5[3][12] } = L4[3][12] + L4[3+1][12] + L4[3+2][12];

assign { L5[0][13+1], L5[2][13] } = L4[0][13] + L4[0+1][13] + L4[0+2][13];
assign { L5[1][13+1], L5[3][13] } = L4[3][13] + L4[3+1][13] + L4[3+2][13];

assign { L5[0][14+1], L5[2][14] } = L4[0][14] + L4[0+1][14] + L4[0+2][14];
assign { L5[1][14+1], L5[3][14] } = L4[3][14] + L4[3+1][14] + L4[3+2][14];

assign { L5[0][15+1], L5[2][15] } = L4[0][15] + L4[0+1][15] + L4[0+2][15];
assign { L5[1][15+1], L5[3][15] } = L4[3][15] + L4[3+1][15] + L4[3+2][15];

assign { L5[0][16+1], L5[2][16] } = L4[0][16] + L4[0+1][16] + L4[0+2][16];
assign { L5[1][16+1], L5[3][16] } = L4[3][16] + L4[3+1][16] + L4[3+2][16];

assign { L5[0][17+1], L5[2][17] } = L4[0][17] + L4[0+1][17] + L4[0+2][17];
assign { L5[1][17+1], L5[3][17] } = L4[3][17] + L4[3+1][17] + L4[3+2][17];

assign { L5[0][18+1], L5[2][18] } = L4[0][18] + L4[0+1][18] + L4[0+2][18];
assign { L5[1][18+1], L5[3][18] } = L4[3][18] + L4[3+1][18] + L4[3+2][18];

assign { L5[0][19+1], L5[2][19] } = L4[0][19] + L4[0+1][19] + L4[0+2][19];
assign { L5[1][19+1], L5[3][19] } = L4[3][19] + L4[3+1][19] + L4[3+2][19];

assign { L5[0][20+1], L5[2][20] } = L4[0][20] + L4[0+1][20] + L4[0+2][20];
assign { L5[1][20+1], L5[3][20] } = L4[3][20] + L4[3+1][20] + L4[3+2][20];

assign { L5[0][21+1], L5[2][21] } = L4[0][21] + L4[0+1][21] + L4[0+2][21];
assign { L5[1][21+1], L5[3][21] } = L4[3][21] + L4[3+1][21] + L4[3+2][21];

assign { L5[0][22+1], L5[2][22] } = L4[0][22] + L4[0+1][22] + L4[0+2][22];
assign { L5[1][22+1], L5[3][22] } = L4[3][22] + L4[3+1][22] + L4[3+2][22];

assign { L5[0][23+1], L5[2][23] } = L4[0][23] + L4[0+1][23] + L4[0+2][23];
assign { L5[1][23+1], L5[3][23] } = L4[3][23] + L4[3+1][23] + L4[3+2][23];

assign { L5[0][24+1], L5[2][24] } = L4[0][24] + L4[0+1][24] + L4[0+2][24];
assign { L5[1][24+1], L5[3][24] } = L4[3][24] + L4[3+1][24] + L4[3+2][24];

assign { L5[0][25+1], L5[2][25] } = L4[0][25] + L4[0+1][25] + L4[0+2][25];
assign { L5[1][25+1], L5[3][25] } = L4[3][25] + L4[3+1][25] + L4[3+2][25];

assign { L5[0][26+1], L5[2][26] } = L4[0][26] + L4[0+1][26] + L4[0+2][26];
assign { L5[1][26+1], L5[3][26] } = L4[3][26] + L4[3+1][26] + L4[3+2][26];

assign { L5[0][27+1], L5[2][27] } = L4[0][27] + L4[0+1][27] + L4[0+2][27];
assign { L5[1][27+1], L5[3][27] } = L4[3][27] + L4[3+1][27] + L4[3+2][27];

assign { L5[0][28+1], L5[2][28] } = L4[0][28] + L4[0+1][28] + L4[0+2][28];
assign { L5[1][28+1], L5[3][28] } = L4[3][28] + L4[3+1][28] + L4[3+2][28];

assign { L5[0][29+1], L5[2][29] } = L4[0][29] + L4[0+1][29] + L4[0+2][29];
assign { L5[1][29+1], L5[3][29] } = L4[3][29] + L4[3+1][29] + L4[3+2][29];

assign { L5[0][30+1], L5[2][30] } = L4[0][30] + L4[0+1][30] + L4[0+2][30];
assign { L5[1][30+1], L5[3][30] } = L4[3][30] + L4[3+1][30] + L4[3+2][30];

assign { L5[0][31+1], L5[2][31] } = L4[0][31] + L4[0+1][31] + L4[0+2][31];
assign { L5[1][31+1], L5[3][31] } = L4[3][31] + L4[3+1][31] + L4[3+2][31];

assign { L5[0][32+1], L5[2][32] } = L4[0][32] + L4[0+1][32] + L4[0+2][32];
assign { L5[1][32+1], L5[3][32] } = L4[3][32] + L4[3+1][32] + L4[3+2][32];

assign { L5[0][33+1], L5[2][33] } = L4[0][33] + L4[0+1][33] + L4[0+2][33];
assign { L5[1][33+1], L5[3][33] } = L4[3][33] + L4[3+1][33] + L4[3+2][33];

assign { L5[0][34+1], L5[2][34] } = L4[0][34] + L4[0+1][34] + L4[0+2][34];
assign { L5[1][34+1], L5[3][34] } = L4[3][34] + L4[3+1][34] + L4[3+2][34];

assign { L5[0][35+1], L5[2][35] } = L4[0][35] + L4[0+1][35] + L4[0+2][35];
assign { L5[1][35+1], L5[3][35] } = L4[3][35] + L4[3+1][35] + L4[3+2][35];

assign { L5[0][36+1], L5[2][36] } = L4[0][36] + L4[0+1][36] + L4[0+2][36];
assign { L5[1][36+1], L5[3][36] } = L4[3][36] + L4[3+1][36] + L4[3+2][36];

assign { L5[0][37+1], L5[2][37] } = L4[0][37] + L4[0+1][37] + L4[0+2][37];
assign { L5[1][37+1], L5[3][37] } = L4[3][37] + L4[3+1][37] + L4[3+2][37];

assign { L5[0][38+1], L5[2][38] } = L4[0][38] + L4[0+1][38] + L4[0+2][38];
assign { L5[1][38+1], L5[3][38] } = L4[3][38] + L4[3+1][38] + L4[3+2][38];

assign { L5[0][39+1], L5[2][39] } = L4[0][39] + L4[0+1][39] + L4[0+2][39];
assign { L5[1][39+1], L5[3][39] } = L4[3][39] + L4[3+1][39] + L4[3+2][39];

assign { L5[0][40+1], L5[2][40] } = L4[0][40] + L4[0+1][40] + L4[0+2][40];
assign { L5[1][40+1], L5[3][40] } = L4[3][40] + L4[3+1][40] + L4[3+2][40];

assign { L5[0][41+1], L5[2][41] } = L4[0][41] + L4[0+1][41] + L4[0+2][41];
assign { L5[1][41+1], L5[3][41] } = L4[3][41] + L4[3+1][41] + L4[3+2][41];

assign { L5[0][42+1], L5[2][42] } = L4[0][42] + L4[0+1][42] + L4[0+2][42];
assign { L5[1][42+1], L5[3][42] } = L4[3][42] + L4[3+1][42] + L4[3+2][42];

assign { L5[0][43+1], L5[2][43] } = L4[0][43] + L4[0+1][43] + L4[0+2][43];
assign L5[3][43] = L4[3][43];

assign L5[1][44] = L4[0][44];
assign L5[2][44] = L4[1][44];
assign L5[3][44] = L4[2][44];

assign L5[0][45] = L4[0][45];
assign L5[1][45] = L4[1][45];

assign L5[0][46] = L4[0][46];


assign L6[0][0] = L5[0][0];

assign L6[0][1] = L5[0][1];
assign L6[1][1] = L5[1][1];

assign L6[0][2] = L5[0][2];
assign L6[1][2] = L5[1][2];
assign L6[2][2] = L5[2][2];

assign { L6[0][3+1], L6[0][3] } = L5[0][3] + L5[0+1][3];
assign L6[1][3] = L5[2][3];
assign L6[2][3] = L5[3][3];

assign { L6[0][4+1], L6[1][4] } = L5[0][4] + L5[0+1][4] + L5[0+2][4];
assign L6[2][4] = L5[3][4];

assign { L6[0][5+1], L6[1][5] } = L5[0][5] + L5[0+1][5] + L5[0+2][5];
assign L6[2][5] = L5[3][5];

assign { L6[0][6+1], L6[1][6] } = L5[0][6] + L5[0+1][6] + L5[0+2][6];
assign L6[2][6] = L5[3][6];

assign { L6[0][7+1], L6[1][7] } = L5[0][7] + L5[0+1][7] + L5[0+2][7];
assign L6[2][7] = L5[3][7];

assign { L6[0][8+1], L6[1][8] } = L5[0][8] + L5[0+1][8] + L5[0+2][8];
assign L6[2][8] = L5[3][8];

assign { L6[0][9+1], L6[1][9] } = L5[0][9] + L5[0+1][9] + L5[0+2][9];
assign L6[2][9] = L5[3][9];

assign { L6[0][10+1], L6[1][10] } = L5[0][10] + L5[0+1][10] + L5[0+2][10];
assign L6[2][10] = L5[3][10];

assign { L6[0][11+1], L6[1][11] } = L5[0][11] + L5[0+1][11] + L5[0+2][11];
assign L6[2][11] = L5[3][11];

assign { L6[0][12+1], L6[1][12] } = L5[0][12] + L5[0+1][12] + L5[0+2][12];
assign L6[2][12] = L5[3][12];

assign { L6[0][13+1], L6[1][13] } = L5[0][13] + L5[0+1][13] + L5[0+2][13];
assign L6[2][13] = L5[3][13];

assign { L6[0][14+1], L6[1][14] } = L5[0][14] + L5[0+1][14] + L5[0+2][14];
assign L6[2][14] = L5[3][14];

assign { L6[0][15+1], L6[1][15] } = L5[0][15] + L5[0+1][15] + L5[0+2][15];
assign L6[2][15] = L5[3][15];

assign { L6[0][16+1], L6[1][16] } = L5[0][16] + L5[0+1][16] + L5[0+2][16];
assign L6[2][16] = L5[3][16];

assign { L6[0][17+1], L6[1][17] } = L5[0][17] + L5[0+1][17] + L5[0+2][17];
assign L6[2][17] = L5[3][17];

assign { L6[0][18+1], L6[1][18] } = L5[0][18] + L5[0+1][18] + L5[0+2][18];
assign L6[2][18] = L5[3][18];

assign { L6[0][19+1], L6[1][19] } = L5[0][19] + L5[0+1][19] + L5[0+2][19];
assign L6[2][19] = L5[3][19];

assign { L6[0][20+1], L6[1][20] } = L5[0][20] + L5[0+1][20] + L5[0+2][20];
assign L6[2][20] = L5[3][20];

assign { L6[0][21+1], L6[1][21] } = L5[0][21] + L5[0+1][21] + L5[0+2][21];
assign L6[2][21] = L5[3][21];

assign { L6[0][22+1], L6[1][22] } = L5[0][22] + L5[0+1][22] + L5[0+2][22];
assign L6[2][22] = L5[3][22];

assign { L6[0][23+1], L6[1][23] } = L5[0][23] + L5[0+1][23] + L5[0+2][23];
assign L6[2][23] = L5[3][23];

assign { L6[0][24+1], L6[1][24] } = L5[0][24] + L5[0+1][24] + L5[0+2][24];
assign L6[2][24] = L5[3][24];

assign { L6[0][25+1], L6[1][25] } = L5[0][25] + L5[0+1][25] + L5[0+2][25];
assign L6[2][25] = L5[3][25];

assign { L6[0][26+1], L6[1][26] } = L5[0][26] + L5[0+1][26] + L5[0+2][26];
assign L6[2][26] = L5[3][26];

assign { L6[0][27+1], L6[1][27] } = L5[0][27] + L5[0+1][27] + L5[0+2][27];
assign L6[2][27] = L5[3][27];

assign { L6[0][28+1], L6[1][28] } = L5[0][28] + L5[0+1][28] + L5[0+2][28];
assign L6[2][28] = L5[3][28];

assign { L6[0][29+1], L6[1][29] } = L5[0][29] + L5[0+1][29] + L5[0+2][29];
assign L6[2][29] = L5[3][29];

assign { L6[0][30+1], L6[1][30] } = L5[0][30] + L5[0+1][30] + L5[0+2][30];
assign L6[2][30] = L5[3][30];

assign { L6[0][31+1], L6[1][31] } = L5[0][31] + L5[0+1][31] + L5[0+2][31];
assign L6[2][31] = L5[3][31];

assign { L6[0][32+1], L6[1][32] } = L5[0][32] + L5[0+1][32] + L5[0+2][32];
assign L6[2][32] = L5[3][32];

assign { L6[0][33+1], L6[1][33] } = L5[0][33] + L5[0+1][33] + L5[0+2][33];
assign L6[2][33] = L5[3][33];

assign { L6[0][34+1], L6[1][34] } = L5[0][34] + L5[0+1][34] + L5[0+2][34];
assign L6[2][34] = L5[3][34];

assign { L6[0][35+1], L6[1][35] } = L5[0][35] + L5[0+1][35] + L5[0+2][35];
assign L6[2][35] = L5[3][35];

assign { L6[0][36+1], L6[1][36] } = L5[0][36] + L5[0+1][36] + L5[0+2][36];
assign L6[2][36] = L5[3][36];

assign { L6[0][37+1], L6[1][37] } = L5[0][37] + L5[0+1][37] + L5[0+2][37];
assign L6[2][37] = L5[3][37];

assign { L6[0][38+1], L6[1][38] } = L5[0][38] + L5[0+1][38] + L5[0+2][38];
assign L6[2][38] = L5[3][38];

assign { L6[0][39+1], L6[1][39] } = L5[0][39] + L5[0+1][39] + L5[0+2][39];
assign L6[2][39] = L5[3][39];

assign { L6[0][40+1], L6[1][40] } = L5[0][40] + L5[0+1][40] + L5[0+2][40];
assign L6[2][40] = L5[3][40];

assign { L6[0][41+1], L6[1][41] } = L5[0][41] + L5[0+1][41] + L5[0+2][41];
assign L6[2][41] = L5[3][41];

assign { L6[0][42+1], L6[1][42] } = L5[0][42] + L5[0+1][42] + L5[0+2][42];
assign L6[2][42] = L5[3][42];

assign { L6[0][43+1], L6[1][43] } = L5[0][43] + L5[0+1][43] + L5[0+2][43];
assign L6[2][43] = L5[3][43];

assign { L6[0][44+1], L6[1][44] } = L5[0][44] + L5[0+1][44] + L5[0+2][44];
assign L6[2][44] = L5[3][44];

assign L6[1][45] = L5[0][45];
assign L6[2][45] = L5[1][45];

assign L6[0][46] = L5[0][46];


assign L7[0][0] = L6[0][0];

assign L7[0][1] = L6[0][1];
assign L7[1][1] = L6[1][1];

assign { L7[0][2+1], L7[0][2] } = L6[0][2] + L6[0+1][2];
assign L7[1][2] = L6[2][2];

assign { L7[0][3+1], L7[1][3] } = L6[0][3] + L6[0+1][3] + L6[0+2][3];

assign { L7[0][4+1], L7[1][4] } = L6[0][4] + L6[0+1][4] + L6[0+2][4];

assign { L7[0][5+1], L7[1][5] } = L6[0][5] + L6[0+1][5] + L6[0+2][5];

assign { L7[0][6+1], L7[1][6] } = L6[0][6] + L6[0+1][6] + L6[0+2][6];

assign { L7[0][7+1], L7[1][7] } = L6[0][7] + L6[0+1][7] + L6[0+2][7];

assign { L7[0][8+1], L7[1][8] } = L6[0][8] + L6[0+1][8] + L6[0+2][8];

assign { L7[0][9+1], L7[1][9] } = L6[0][9] + L6[0+1][9] + L6[0+2][9];

assign { L7[0][10+1], L7[1][10] } = L6[0][10] + L6[0+1][10] + L6[0+2][10];

assign { L7[0][11+1], L7[1][11] } = L6[0][11] + L6[0+1][11] + L6[0+2][11];

assign { L7[0][12+1], L7[1][12] } = L6[0][12] + L6[0+1][12] + L6[0+2][12];

assign { L7[0][13+1], L7[1][13] } = L6[0][13] + L6[0+1][13] + L6[0+2][13];

assign { L7[0][14+1], L7[1][14] } = L6[0][14] + L6[0+1][14] + L6[0+2][14];

assign { L7[0][15+1], L7[1][15] } = L6[0][15] + L6[0+1][15] + L6[0+2][15];

assign { L7[0][16+1], L7[1][16] } = L6[0][16] + L6[0+1][16] + L6[0+2][16];

assign { L7[0][17+1], L7[1][17] } = L6[0][17] + L6[0+1][17] + L6[0+2][17];

assign { L7[0][18+1], L7[1][18] } = L6[0][18] + L6[0+1][18] + L6[0+2][18];

assign { L7[0][19+1], L7[1][19] } = L6[0][19] + L6[0+1][19] + L6[0+2][19];

assign { L7[0][20+1], L7[1][20] } = L6[0][20] + L6[0+1][20] + L6[0+2][20];

assign { L7[0][21+1], L7[1][21] } = L6[0][21] + L6[0+1][21] + L6[0+2][21];

assign { L7[0][22+1], L7[1][22] } = L6[0][22] + L6[0+1][22] + L6[0+2][22];

assign { L7[0][23+1], L7[1][23] } = L6[0][23] + L6[0+1][23] + L6[0+2][23];

assign { L7[0][24+1], L7[1][24] } = L6[0][24] + L6[0+1][24] + L6[0+2][24];

assign { L7[0][25+1], L7[1][25] } = L6[0][25] + L6[0+1][25] + L6[0+2][25];

assign { L7[0][26+1], L7[1][26] } = L6[0][26] + L6[0+1][26] + L6[0+2][26];

assign { L7[0][27+1], L7[1][27] } = L6[0][27] + L6[0+1][27] + L6[0+2][27];

assign { L7[0][28+1], L7[1][28] } = L6[0][28] + L6[0+1][28] + L6[0+2][28];

assign { L7[0][29+1], L7[1][29] } = L6[0][29] + L6[0+1][29] + L6[0+2][29];

assign { L7[0][30+1], L7[1][30] } = L6[0][30] + L6[0+1][30] + L6[0+2][30];

assign { L7[0][31+1], L7[1][31] } = L6[0][31] + L6[0+1][31] + L6[0+2][31];

assign { L7[0][32+1], L7[1][32] } = L6[0][32] + L6[0+1][32] + L6[0+2][32];

assign { L7[0][33+1], L7[1][33] } = L6[0][33] + L6[0+1][33] + L6[0+2][33];

assign { L7[0][34+1], L7[1][34] } = L6[0][34] + L6[0+1][34] + L6[0+2][34];

assign { L7[0][35+1], L7[1][35] } = L6[0][35] + L6[0+1][35] + L6[0+2][35];

assign { L7[0][36+1], L7[1][36] } = L6[0][36] + L6[0+1][36] + L6[0+2][36];

assign { L7[0][37+1], L7[1][37] } = L6[0][37] + L6[0+1][37] + L6[0+2][37];

assign { L7[0][38+1], L7[1][38] } = L6[0][38] + L6[0+1][38] + L6[0+2][38];

assign { L7[0][39+1], L7[1][39] } = L6[0][39] + L6[0+1][39] + L6[0+2][39];

assign { L7[0][40+1], L7[1][40] } = L6[0][40] + L6[0+1][40] + L6[0+2][40];

assign { L7[0][41+1], L7[1][41] } = L6[0][41] + L6[0+1][41] + L6[0+2][41];

assign { L7[0][42+1], L7[1][42] } = L6[0][42] + L6[0+1][42] + L6[0+2][42];

assign { L7[0][43+1], L7[1][43] } = L6[0][43] + L6[0+1][43] + L6[0+2][43];

assign { L7[0][44+1], L7[1][44] } = L6[0][44] + L6[0+1][44] + L6[0+2][44];

assign { L7[0][45+1], L7[1][45] } = L6[0][45] + L6[0+1][45] + L6[0+2][45];

assign L7[1][46] = L6[0][46];

endmodule
