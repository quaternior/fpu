module FMUL_add(
    
);

endmodule